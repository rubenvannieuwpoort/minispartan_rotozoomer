----------------------------------------------------------------------------------
-- Engineer:   Ruben van Nieuwpoort <benoncoffee@gmail.com>
-- 
-- Module Name: lut - Behavioral 
-- Description: A lookup table for the sine and cosine at 1024 angles.
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity lut is
	generic (
		frac_bits  : natural;
		lut_size  : natural
	);
	port(
		angle : in  unsigned( 8 downto 0);
		sin   : out signed(15 downto 0);
		cos   : out signed(15 downto 0)
	);
end lut;

architecture Behavioral of lut is
	
	constant int_bits : natural := 2;
	constant total_bits : natural := int_bits + frac_bits;

	type memory is array(0 to lut_size - 1) of std_logic_vector(2 * total_bits - 1 downto 0);
	signal rom : memory := 
	(
		"00000000000000000100000000000000", "00000000110010010011111111111110", "00000001100100100011111111111011", "00000010010110110011111111110100",
		"00000011001000110011111111101100", "00000011111011000011111111100001", "00000100101101010011111111010011", "00000101011111010011111111000011",
		"00000110010001010011111110110001", "00000111000011010011111110011100", "00000111110101010011111110000100", "00001000100111000011111101101010",
		"00001001011001000011111101001110", "00001010001010100011111100101111", "00001010111100010011111100001110", "00001011101101100011111011101011",
		"00001100011111000011111011000101", "00001101010000010011111010011100", "00001110000001010011111001110001", "00001110110010010011111001000100",
		"00001111100011000011111000010100", "00010000010011110011110111100010", "00010001000100010011110110101110", "00010001110100110011110101110111",
		"00010010100101000011110100111110", "00010011010101000011110100000010", "00010100000100110011110011000101", "00010100110100010011110010000100",
		"00010101100011110011110001000010", "00010110010011000011101111111101", "00010111000010000011101110110110", "00010111110000110011101101101100",
		"00011000011111010011101100100000", "00011001001101110011101011010010", "00011001111011110011101010000010", "00011010101001100011101000101111",
		"00011011010111010011100111011010", "00011100000100100011100110000011", "00011100110001100011100100101010", "00011101011110010011100011001111",
		"00011110001010110011100001110001", "00011110110111000011100000010001", "00011111100010110011011110101111", "00100000001110010011011101001011",
		"00100000111001110011011011100101", "00100001100100100011011001111100", "00100010001111010011011000010010", "00100010111001100011010110100101",
		"00100011100011100011010100110110", "00100100001101000011010011000110", "00100100110110100011010001010011", "00100101011111010011001111011110",
		"00100110000111110011001101100111", "00100110110000000011001011101110", "00100111010111110011001001110100", "00100111111111010011000111110111",
		"00101000100110010011000101111001", "00101001001101000011000011111000", "00101001110011010011000001110110", "00101010011001010010111111110001",
		"00101010111110100010111101101011", "00101011100011100010111011100011", "00101100001000010010111001011010", "00101100101100100010110111001110",
		"00101101010000010010110101000001", "00101101110011100010110010110010", "00101110010110100010110000100001", "00101110111000110010101110001110",
		"00101111011010110010101011111010", "00101111111100010010101001100101", "00110000011101100010100111001101", "00110000111110000010100100110100",
		"00110001011110010010100010011001", "00110001111101110010011111111101", "00110010011101000010011101011111", "00110010111011100010011011000000",
		"00110011011001110010011000011111", "00110011110111100010010101111101", "00110100010100110010010011011010", "00110100110001100010010000110100",
		"00110101001101100010001110001110", "00110101101001010010001011100110", "00110110000100100010001000111101", "00110110011111000010000110010010",
		"00110110111001010010000011100111", "00110111010010110010000000111001", "00110111101011110001111110001011", "00111000000100010001111011011100",
		"00111000011100010001111000101011", "00111000110011110001110101111001", "00111001001010100001110011000110", "00111001100000110001110000010010",
		"00111001110110100001101101011101", "00111010001011110001101010100110", "00111010100000100001100111101111", "00111010110100100001100100110111",
		"00111011001000000001100001111101", "00111011011011000001011111000011", "00111011101101100001011100001000", "00111011111111010001011001001100",
		"00111100010000100001010110001111", "00111100100001000001010011010001", "00111100110001010001010000010011", "00111101000000100001001101010100",
		"00111101001111100001001010010100", "00111101011101110001000111010011", "00111101101011100001000100010001", "00111101111000100001000001001111",
		"00111110000101000000111110001100", "00111110010001000000111011001001", "00111110011100010000111000000101", "00111110100111000000110101000001",
		"00111110110001010000110001111100", "00111110111010110000101110110110", "00111111000011100000101011110001", "00111111001011110000101000101010",
		"00111111010011100000100101100100", "00111111011010100000100010011100", "00111111100001000000011111010101", "00111111100111000000011100001101",
		"00111111101100010000011001000101", "00111111110000110000010101111101", "00111111110100110000010010110101", "00111111111000010000001111101100",
		"00111111111011000000001100100011", "00111111111101000000001001011011", "00111111111110110000000110010010", "00111111111111100000000011001001",
		"01000000000000000000000000000000", "00111111111111101111111100110111", "00111111111110111111111001101110", "00111111111101001111110110100101",
		"00111111111011001111110011011101", "00111111111000011111110000010100", "00111111110100111111101101001011", "00111111110000111111101010000011",
		"00111111101100011111100110111011", "00111111100111001111100011110011", "00111111100001001111100000101011", "00111111011010101111011101100100",
		"00111111010011101111011010011100", "00111111001011111111010111010110", "00111111000011101111010100001111", "00111110111010111111010001001010",
		"00111110110001011111001110000100", "00111110100111001111001010111111", "00111110011100011111000111111011", "00111110010001001111000100110111",
		"00111110000101001111000001110100", "00111101111000101110111110110001", "00111101101011101110111011101111", "00111101011101111110111000101101",
		"00111101001111101110110101101100", "00111101000000101110110010101100", "00111100110001011110101111101101", "00111100100001001110101100101111",
		"00111100010000101110101001110001", "00111011111111011110100110110100", "00111011101101101110100011111000", "00111011011011001110100000111101",
		"00111011001000001110011110000011", "00111010110100101110011011001001", "00111010100000101110011000010001", "00111010001011111110010101011010",
		"00111001110110101110010010100011", "00111001100000111110001111101110", "00111001001010101110001100111010", "00111000110011111110001010000111",
		"00111000011100011110000111010101", "00111000000100011110000100100100", "00110111101011111110000001110101", "00110111010010111101111111000111",
		"00110110111001011101111100011001", "00110110011111001101111001101110", "00110110000100101101110111000011", "00110101101001011101110100011010",
		"00110101001101101101110001110010", "00110100110001101101101111001100", "00110100010100111101101100100110", "00110011110111101101101010000011",
		"00110011011001111101100111100001", "00110010111011101101100101000000", "00110010011101001101100010100001", "00110001111101111101100000000011",
		"00110001011110011101011101100111", "00110000111110001101011011001100", "00110000011101101101011000110011", "00101111111100011101010110011011",
		"00101111011010111101010100000110", "00101110111000111101010001110010", "00101110010110101101001111011111", "00101101110011101101001101001110",
		"00101101010000011101001010111111", "00101100101100101101001000110010", "00101100001000011101000110100110", "00101011100011101101000100011101",
		"00101010111110101101000010010101", "00101010011001011101000000001111", "00101001110011011100111110001010", "00101001001101001100111100001000",
		"00101000100110011100111010000111", "00100111111111011100111000001001", "00100111010111111100110110001100", "00100110110000001100110100010010",
		"00100110000111111100110010011001", "00100101011111011100110000100010", "00100100110110101100101110101101", "00100100001101001100101100111010",
		"00100011100011101100101011001010", "00100010111001101100101001011011", "00100010001111011100100111101110", "00100001100100101100100110000100",
		"00100000111001111100100100011011", "00100000001110011100100010110101", "00011111100010111100100001010001", "00011110110111001100011111101111",
		"00011110001010111100011110001111", "00011101011110011100011100110001", "00011100110001101100011011010110", "00011100000100101100011001111101",
		"00011011010111011100011000100110", "00011010101001101100010111010001", "00011001111011111100010101111110", "00011001001101111100010100101110",
		"00011000011111011100010011100000", "00010111110000111100010010010100", "00010111000010001100010001001010", "00010110010011001100010000000011",
		"00010101100011111100001110111110", "00010100110100011100001101111100", "00010100000100111100001100111011", "00010011010101001100001011111110",
		"00010010100101001100001011000010", "00010001110100111100001010001001", "00010001000100011100001001010010", "00010000010011111100001000011110",
		"00001111100011001100000111101100", "00001110110010011100000110111100", "00001110000001011100000110001111", "00001101010000011100000101100100",
		"00001100011111001100000100111011", "00001011101101101100000100010101", "00001010111100011100000011110010", "00001010001010101100000011010001",
		"00001001011001001100000010110010", "00001000100111001100000010010110", "00000111110101011100000001111100", "00000111000011011100000001100100",
		"00000110010001011100000001001111", "00000101011111011100000000111101", "00000100101101011100000000101101", "00000011111011001100000000011111",
		"00000011001000111100000000010100", "00000010010110111100000000001100", "00000001100100101100000000000101", "00000000110010011100000000000010",
		"00000000000000001100000000000000", "11111111001101111100000000000010", "11111110011011101100000000000101", "11111101101001011100000000001100",
		"11111100110111011100000000010100", "11111100000101001100000000011111", "11111011010010111100000000101101", "11111010100000111100000000111101",
		"11111001101110111100000001001111", "11111000111100111100000001100100", "11111000001010111100000001111100", "11110111011001001100000010010110",
		"11110110100111001100000010110010", "11110101110101101100000011010001", "11110101000011111100000011110010", "11110100010010101100000100010101",
		"11110011100001001100000100111011", "11110010101111111100000101100100", "11110001111110111100000110001111", "11110001001101111100000110111100",
		"11110000011101001100000111101100", "11101111101100011100001000011110", "11101110111011111100001001010010", "11101110001011011100001010001001",
		"11101101011011001100001011000010", "11101100101011001100001011111110", "11101011111011011100001100111011", "11101011001011111100001101111100",
		"11101010011100011100001110111110", "11101001101101001100010000000011", "11101000111110001100010001001010", "11101000001111011100010010010100",
		"11100111100000111100010011100000", "11100110110010011100010100101110", "11100110000100011100010101111110", "11100101010110101100010111010001",
		"11100100101000111100011000100110", "11100011111011101100011001111101", "11100011001110101100011011010110", "11100010100001111100011100110001",
		"11100001110101011100011110001111", "11100001001001001100011111101111", "11100000011101011100100001010001", "11011111110001111100100010110101",
		"11011111000110011100100100011011", "11011110011011101100100110000100", "11011101110000111100100111101110", "11011101000110101100101001011011",
		"11011100011100101100101011001010", "11011011110011001100101100111010", "11011011001001101100101110101101", "11011010100000111100110000100010",
		"11011001111000011100110010011001", "11011001010000001100110100010010", "11011000101000011100110110001100", "11011000000000111100111000001001",
		"11010111011001111100111010000111", "11010110110011001100111100001000", "11010110001100111100111110001010", "11010101100110111101000000001111",
		"11010101000001101101000010010101", "11010100011100101101000100011101", "11010011110111111101000110100110", "11010011010011101101001000110010",
		"11010010101111111101001010111111", "11010010001100101101001101001110", "11010001101001101101001111011111", "11010001000111011101010001110010",
		"11010000100101011101010100000110", "11010000000011111101010110011011", "11001111100010101101011000110011", "11001111000010001101011011001100",
		"11001110100001111101011101100111", "11001110000010011101100000000011", "11001101100011001101100010100001", "11001101000100101101100101000000",
		"11001100100110011101100111100001", "11001100001000101101101010000011", "11001011101011011101101100100110", "11001011001110101101101111001100",
		"11001010110010101101110001110010", "11001010010110111101110100011010", "11001001111011101101110111000011", "11001001100001001101111001101110",
		"11001001000110111101111100011001", "11001000101101011101111111000111", "11001000010100011110000001110101", "11000111111011111110000100100100",
		"11000111100011111110000111010101", "11000111001100011110001010000111", "11000110110101101110001100111010", "11000110011111011110001111101110",
		"11000110001001101110010010100011", "11000101110100011110010101011010", "11000101011111101110011000010001", "11000101001011101110011011001001",
		"11000100111000001110011110000011", "11000100100101001110100000111101", "11000100010010101110100011111000", "11000100000000111110100110110100",
		"11000011101111101110101001110001", "11000011011111001110101100101111", "11000011001110111110101111101101", "11000010111111101110110010101100",
		"11000010110000101110110101101100", "11000010100010011110111000101101", "11000010010100101110111011101111", "11000010000111101110111110110001",
		"11000001111011001111000001110100", "11000001101111001111000100110111", "11000001100011111111000111111011", "11000001011001001111001010111111",
		"11000001001110111111001110000100", "11000001000101011111010001001010", "11000000111100101111010100001111", "11000000110100011111010111010110",
		"11000000101100101111011010011100", "11000000100101101111011101100100", "11000000011111001111100000101011", "11000000011001001111100011110011",
		"11000000010011111111100110111011", "11000000001111011111101010000011", "11000000001011011111101101001011", "11000000000111111111110000010100",
		"11000000000101001111110011011101", "11000000000011001111110110100101", "11000000000001011111111001101110", "11000000000000101111111100110111",
		"11000000000000000000000000000000", "11000000000000100000000011001001", "11000000000001010000000110010010", "11000000000011000000001001011011",
		"11000000000101000000001100100011", "11000000000111110000001111101100", "11000000001011010000010010110101", "11000000001111010000010101111101",
		"11000000010011110000011001000101", "11000000011001000000011100001101", "11000000011111000000011111010101", "11000000100101100000100010011100",
		"11000000101100100000100101100100", "11000000110100010000101000101010", "11000000111100100000101011110001", "11000001000101010000101110110110",
		"11000001001110110000110001111100", "11000001011001000000110101000001", "11000001100011110000111000000101", "11000001101111000000111011001001",
		"11000001111011000000111110001100", "11000010000111100001000001001111", "11000010010100100001000100010001", "11000010100010010001000111010011",
		"11000010110000100001001010010100", "11000010111111100001001101010100", "11000011001110110001010000010011", "11000011011111000001010011010001",
		"11000011101111100001010110001111", "11000100000000110001011001001100", "11000100010010100001011100001000", "11000100100101000001011111000011",
		"11000100111000000001100001111101", "11000101001011100001100100110111", "11000101011111100001100111101111", "11000101110100010001101010100110",
		"11000110001001100001101101011101", "11000110011111010001110000010010", "11000110110101100001110011000110", "11000111001100010001110101111001",
		"11000111100011110001111000101011", "11000111111011110001111011011100", "11001000010100010001111110001011", "11001000101101010010000000111001",
		"11001001000110110010000011100111", "11001001100001000010000110010010", "11001001111011100010001000111101", "11001010010110110010001011100110",
		"11001010110010100010001110001110", "11001011001110100010010000110100", "11001011101011010010010011011010", "11001100001000100010010101111101",
		"11001100100110010010011000011111", "11001101000100100010011011000000", "11001101100011000010011101011111", "11001110000010010010011111111101",
		"11001110100001110010100010011001", "11001111000010000010100100110100", "11001111100010100010100111001101", "11010000000011110010101001100101",
		"11010000100101010010101011111010", "11010001000111010010101110001110", "11010001101001100010110000100001", "11010010001100100010110010110010",
		"11010010101111110010110101000001", "11010011010011100010110111001110", "11010011110111110010111001011010", "11010100011100100010111011100011",
		"11010101000001100010111101101011", "11010101100110110010111111110001", "11010110001100110011000001110110", "11010110110011000011000011111000",
		"11010111011001110011000101111001", "11011000000000110011000111110111", "11011000101000010011001001110100", "11011001010000000011001011101110",
		"11011001111000010011001101100111", "11011010100000110011001111011110", "11011011001001100011010001010011", "11011011110011000011010011000110",
		"11011100011100100011010100110110", "11011101000110100011010110100101", "11011101110000110011011000010010", "11011110011011100011011001111100",
		"11011111000110010011011011100101", "11011111110001110011011101001011", "11100000011101010011011110101111", "11100001001001000011100000010001",
		"11100001110101010011100001110001", "11100010100001110011100011001111", "11100011001110100011100100101010", "11100011111011100011100110000011",
		"11100100101000110011100111011010", "11100101010110100011101000101111", "11100110000100010011101010000010", "11100110110010010011101011010010",
		"11100111100000110011101100100000", "11101000001111010011101101101100", "11101000111110000011101110110110", "11101001101101000011101111111101",
		"11101010011100010011110001000010", "11101011001011110011110010000100", "11101011111011010011110011000101", "11101100101011000011110100000010",
		"11101101011011000011110100111110", "11101110001011010011110101110111", "11101110111011110011110110101110", "11101111101100010011110111100010",
		"11110000011101000011111000010100", "11110001001101110011111001000100", "11110001111110110011111001110001", "11110010101111110011111010011100",
		"11110011100001000011111011000101", "11110100010010100011111011101011", "11110101000011110011111100001110", "11110101110101100011111100101111",
		"11110110100111000011111101001110", "11110111011001000011111101101010", "11111000001010110011111110000100", "11111000111100110011111110011100",
		"11111001101110110011111110110001", "11111010100000110011111111000011", "11111011010010110011111111010011", "11111100000101000011111111100001",
		"11111100110111010011111111101100", "11111101101001010011111111110100", "11111110011011100011111111111011", "11111111001101110011111111111110"
	);
begin
	sin <= signed(rom(to_integer(unsigned(angle)))(2 * total_bits - 1 downto total_bits));
	cos <= signed(rom(to_integer(unsigned(angle)))(total_bits - 1 downto 0));
end Behavioral;

