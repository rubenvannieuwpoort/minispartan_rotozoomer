----------------------------------------------------------------------------------
-- Engineer:   Ruben van Nieuwpoort <benoncoffee@gmail.com>
-- 
-- Module Name: texture_uv_lut - Behavioral 
-- Description: A lookup table for the U and V values of the famous Lena picture.
----------------------------------------------------------------------------------

library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity texture_uv_lut is
	port(
		clk : std_logic;
		address : in std_logic_vector(13 downto 0);
		data : out std_logic_vector(15 downto 0)
	);
end texture_uv_lut;

architecture Behavioral of texture_uv_lut is
	type memory is array(0 to 16383) of std_logic_vector(15 downto 0);
	signal rom : memory := 
	(
		"1010010001111101", "1010001101111101", "1010001001111110", "1010001001111110", "1010001001111110", "1010001001111110", "1010001101111101", "1010001001111110", "1010001001111110", "1010001101111110", "1010001101111101", "1010010001111101", "1010010001111101", "1010001101111110", "1010001101111111", "1010001101111111", "1010001101111110", "1010001001111110", "1001111001111101", "1001100101111101", "1001011101111101", "1001011101111101", "1001100001111101", "1001100001111101", "1001100001111101", "1001100001111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1010000101111101", "1010000101111101", "1010010001111101", "1010010101111101", "1010011001111101", "1010011101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010010001111110", "1010010001111101", "1010010001111101", "1010001101111111", "1010010001111101", "1010010101111101", "1010010101111110", "1010001010000000", "1001111010000101", "1001100110000101", "1001100110000100", "1001111010000100", "1010000101111111", "1001110001111110", "1001110001111110", "1001110001111101", "1001101101111110", "1001101001111110", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111110", "1001110001111101", "1001111001111101", "1001111101111101", "1001111001111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111101111101", "1001111101111111", "1001101110000001", "1001100110000001", "1001110001111111", "1001010001111111", "1010010001111101", "1010001101111101", "1010001001111110", "1010001001111110", "1010001001111110", "1010001001111110", "1010001001111110", "1010001001111110", "1010001001111110", "1010001001111110", "1010001101111101", "1010010001111101", "1010001101111101", "1010010001111101", "1010001101111111", "1010010001111101", "1010001001111110", "1010000001111110", "1001101101111110", "1001011101111101", "1001100001111101", "1001100001111101", "1001100001111101", "1001100001111101", "1001100001111101", "1001100101111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000001111101", "1001111101111101", "1010000001111101", "1010000001111101", "1001111101111101", "1010000001111101", "1001111101111101", "1010000001111101", "1001111101111101", "1010000001111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001111101111101", "1010001001111101", "1010001101111101", "1010010001111101", "1010010101111101", "1010011001111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010010001111110", "1010010001111110", "1010010001111110", "1010010001111110", "1010010101111101", "1010010101111101", "1010010101111111", "1010000110000001", "1001110110000100", "1001101010000100", "1001101010000100", "1001111110000001", "1001111001111111", "1001110001111110", "1001110001111101", "1001110001111110", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111110", "1001111001111101", "1001111001111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001111001111101", "1010000001111101", "1001111001111111", "1001100110000001", "1001101010000000", "1001110001111111", "1010001101111101", "1010001001111110", "1010001001111110", "1010001001111110", "1010001001111110", "1010001101111101", "1010001101111101", "1010001001111110", "1010001001111110", "1010001001111110", "1010001101111101", "1010001101111101", "1010001101111110", "1010001101111111", "1010010001111110", "1010001101111110", "1010000101111110", "1001110101111101", "1001100001111101", "1001100001111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000101111101", "1010000001111101", "1010000101111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000001111101", "1001111101111101", "1001111101111101", "1010000101111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000001111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110001111101", "1001110101111101", "1010000001111101", "1010001001111101", "1010010001111101", "1010010101111101", "1010010101111110", "1010011001111101", "1010010101111110", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010010101111101", "1010010001111110", "1010001101111110", "1010010101111101", "1010010001111110", "1010010001111101", "1010010101111101", "1010010101111110", "1010010001111111", "1001111110000100", "1001110010000101", "1001101010000101", "1001110110000100", "1001111101111111", "1001111001111110", "1001110101111110", "1001110001111110", "1001110001111110", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111001111101", "1001110001111110", "1001110101111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001111101111101", "1010000001111111", "1001110010000000", "1001100110000001", "1001101101111111", "1010001001111110", "1010001101111110", "1010001101111101", "1010001001111110", "1010001101111110", "1010001101111101", "1010001001111110", "1010001001111110", "1010001001111110", "1010001101111101", "1010001001111110", "1010001101111101", "1010001101111110", "1010001101111111", "1010001101111111", "1010001101111110", "1001111101111110", "1001100101111101", "1001011101111101", "1001100101111101", "1001101001111101", "1001101001111101", "1001100101111101", "1001101101111100", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010001001111100", "1010001001111101", "1010001001111100", "1010001101111101", "1010001001111101", "1010000101111101", "1010001001111101", "1010001001111101", "1010001101111100", "1010001101111101", "1010001101111100", "1010001001111101", "1010001001111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000001111101", "1010000001111101", "1001111101111110", "1010000001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110001111101", "1001111101111101", "1010001001111101", "1010010001111101", "1010010001111101", "1010010101111101", "1010011001111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010101111101", "1010010001111101", "1010010001111110", "1010010001111110", "1010010001111101", "1010010001111110", "1010010001111110", "1010010001111101", "1010010001111110", "1010010101111111", "1010001110000001", "1001111010000100", "1001101010000101", "1001101010000101", "1001111010000011", "1001111101111111", "1001110101111111", "1001110001111110", "1001110001111110", "1001110001111101", "1001110001111110", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001110101111110", "1001111001111101", "1001110101111101", "1001110001111110", "1001110001111101", "1001111101111100", "1001111001111101", "1001110101111101", "1001111101111101", "1001111101111110", "1001111101111111", "1001101010000001", "1001100110000001", "1010001101111101", "1010001001111110", "1010001001111110", "1010001001111110", "1010001101111101", "1010001101111101", "1010001101111101", "1010001001111110", "1010001001111110", "1010001101111101", "1010001101111101", "1010001101111110", "1010001101111111", "1010010001111111", "1010010001111110", "1010001101111110", "1001111001111101", "1001011101111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000101111101", "1010000101111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010001001111100", "1010001001111100", "1010001001111101", "1010001101111100", "1010001101111100", "1010001001111101", "1010001101111101", "1010001001111101", "1010010001111100", "1010001101111100", "1010010001111100", "1010001001111101", "1010001001111101", "1010001001111100", "1010001001111101", "1010001001111100", "1010000101111101", "1010000101111101", "1010000101111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010001001111100", "1010001001111100", "1010001001111101", "1010001001111100", "1010001001111101", "1010001001111100", "1010000101111101", "1010000101111101", "1010000001111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001111101111101", "1010001001111101", "1010010001111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111110", "1010010101111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010010001111110", "1010010001111111", "1010010101111111", "1010000110000011", "1001110010000110", "1001100110000110", "1001100110000100", "1001111110000000", "1001111001111111", "1001110101111110", "1001110001111110", "1001110001111110", "1001110001111110", "1001110101111101", "1001110101111110", "1001110001111110", "1001110001111110", "1001110001111110", "1001111001111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001110101111110", "1001110101111101", "1001111101111101", "1001111001111101", "1001111001111101", "1001111101111111", "1001110001111111", "1001100110000001", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001001111110", "1010001001111110", "1010001001111110", "1010001001111110", "1010001101111101", "1010001101111111", "1010010001111111", "1010010001111111", "1010010001111110", "1010001001111110", "1001110001111101", "1001011101111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001101101111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000101111100", "1010000101111101", "1010000101111101", "1010001001111101", "1010000101111101", "1010001101111100", "1010001101111100", "1010001101111011", "1010001101111100", "1010001101111011", "1010001101111100", "1010001101111100", "1010001101111100", "1010010001111100", "1010010001111011", "1010001101111100", "1010001001111101", "1010001001111100", "1010001101111100", "1010001001111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010001001111100", "1010001001111100", "1010001001111100", "1010000101111101", "1010001001111101", "1010000101111101", "1010000001111101", "1010000001111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1010000101111101", "1010001001111101", "1010010001111101", "1010010001111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010101111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010010001111110", "1010010001111110", "1010001110000000", "1001111010000100", "1001100110000101", "1001011110000101", "1001110010000100", "1001111101111111", "1001111001111110", "1001110101111110", "1001110101111110", "1001110101111110", "1001110101111110", "1001110101111110", "1001110101111101", "1001110001111110", "1001110001111110", "1001110101111110", "1001110101111110", "1001111001111101", "1001110101111110", "1001110101111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111001111101", "1001111101111101", "1001111101111111", "1001101110000000", "1010001101111110", "1010001101111101", "1010001001111110", "1010001101111101", "1010001101111101", "1010001101111101", "1010001001111101", "1010001001111110", "1010001001111110", "1010001101111101", "1010001001111111", "1010010001111111", "1010010001111111", "1010010001111111", "1010010001111110", "1010000101111110", "1001110001111101", "1001100001111101", "1001100001111101", "1001100101111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000101111101", "1010000101111101", "1010000101111100", "1010000101111101", "1010001001111100", "1010000101111100", "1010001001111101", "1010001101111100", "1010001101111100", "1010001101111100", "1010001101111100", "1010010001111011", "1010001101111100", "1010010001111100", "1010001101111100", "1010010001111100", "1010010001111100", "1010010001111100", "1010010001111100", "1010001001111100", "1010001101111100", "1010001001111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111100", "1010001001111100", "1010001001111100", "1010001001111100", "1010010001111011", "1010001001111100", "1010001001111101", "1010001001111100", "1010000101111101", "1010000101111101", "1010000001111101", "1010000101111101", "1010000001111101", "1010000001111101", "1001111101111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001110001111100", "1001110001111101", "1001111101111101", "1010000101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010101111110", "1010010101111110", "1010010101111101", "1010011001111101", "1010010101111101", "1010010001111101", "1010010001111110", "1010010001111110", "1010010001111110", "1010010001111111", "1010000110000001", "1001110010000101", "1001100010000101", "1001100110000101", "1001111110000010", "1001111101111111", "1001110101111111", "1001110101111110", "1001111001111110", "1001111001111101", "1001110101111101", "1001110101111110", "1001110001111101", "1001110001111110", "1001111001111101", "1001111001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001100001111111", "1010001101111101", "1010001001111110", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001001111110", "1010001001111110", "1010001101111110", "1010001101111111", "1010001101111111", "1010010001111111", "1010010001111111", "1010010001111111", "1010000101111101", "1001110001111101", "1001100001111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111100", "1001110001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010001001111100", "1010001001111100", "1010001001111100", "1010001001111100", "1010001001111100", "1010001101111100", "1010010001111011", "1010010001111100", "1010010001111011", "1010010001111011", "1010010001111011", "1010001101111011", "1010010001111100", "1010010001111100", "1010010001111100", "1010010001111011", "1010001101111100", "1010001101111100", "1010001001111100", "1010001001111100", "1010001001111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111100", "1010001001111101", "1010001001111100", "1010001001111100", "1010001101111100", "1010001001111101", "1010001001111100", "1010001001111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111100", "1001110001111101", "1001110001111101", "1001110101111101", "1010000001111101", "1010000101111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010101111101", "1010011001111101", "1010010101111110", "1010010101111110", "1010010101111110", "1010011001111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111110", "1010001101111111", "1001111110000100", "1001101010000110", "1001100110000101", "1001101110000100", "1010000010000000", "1001111001111111", "1001111001111110", "1001111001111110", "1001110101111110", "1001110101111110", "1001110101111111", "1001110001111110", "1001110101111101", "1001110001111110", "1001111001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001101001111101", "1000111101111111", "1000010001111111", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001001111110", "1010001101111101", "1010001101111111", "1010001101111111", "1010010001111111", "1010001101111111", "1010010001111111", "1010001101111110", "1010000101111110", "1001110001111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000101111101", "1010001001111100", "1010000101111100", "1010001001111101", "1010001101111011", "1010001001111100", "1010010001111011", "1010001101111100", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111100", "1010010001111011", "1010010001111011", "1010001101111100", "1010010001111100", "1010010001111011", "1010010001111011", "1010001101111100", "1010001101111100", "1010001001111100", "1010001001111100", "1010001001111101", "1010000101111101", "1010000101111100", "1010000101111101", "1010000101111101", "1010001001111100", "1010001001111101", "1010001101111011", "1010001101111100", "1010001101111100", "1010001001111101", "1010001101111100", "1010001001111100", "1010001001111100", "1010000101111100", "1010000101111101", "1010000101111101", "1010000001111101", "1010000101111101", "1010000001111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1010000101111101", "1010001101111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111110", "1010011001111110", "1010011001111110", "1010010101111101", "1010011001111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010001101111101", "1010010001111101", "1010001101111110", "1010000110000001", "1001110110000101", "1001100110000101", "1001100010000110", "1001110110000100", "1010000001111111", "1001111001111111", "1001111001111110", "1001111001111110", "1001111001111110", "1001111001111110", "1001111001111101", "1001111001111101", "1001110001111110", "1001110101111101", "1001110101111110", "1001111001111110", "1001111101111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001100101111101", "1000101101111111", "1000000101111111", "0111111101111111", "1010001001111110", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111110", "1010001101111101", "1010001001111110", "1010001001111110", "1010001001111111", "1010001001111111", "1010001001111111", "1010001101111111", "1010010001111110", "1010001101111110", "1010000101111110", "1001110001111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000101111101", "1010000101111101", "1010001001111100", "1010001001111100", "1010001101111011", "1010010001111011", "1010001101111100", "1010001101111011", "1010010001111100", "1010010001111011", "1010010001111011", "1010010001111100", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111100", "1010001101111100", "1010001101111100", "1010001101111100", "1010010001111100", "1010001001111100", "1010001001111100", "1010000101111100", "1010000101111101", "1010001001111100", "1010001001111100", "1010010001111011", "1010001001111100", "1010001101111011", "1010001001111100", "1010010001111011", "1010010001111100", "1010001101111100", "1010001001111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000001111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1010000001111101", "1010000101111101", "1010001101111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010101111110", "1010010101111111", "1010011001111110", "1010011001111101", "1010010101111101", "1010010101111110", "1010010101111110", "1010010101111101", "1010010101111101", "1010010001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111111", "1010000010000011", "1001101010000101", "1001100010000101", "1001100110000101", "1001111110000001", "1001111101111111", "1001110101111111", "1001111001111110", "1001111101111101", "1001110101111110", "1001111001111110", "1001111001111110", "1001110101111110", "1001110101111101", "1001110101111110", "1001111001111110", "1001111101111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001011101111110", "1000100001111111", "1000000101111111", "0111111101111111", "0111111101111111", "1010001001111110", "1010001101111101", "1010001101111101", "1010001101111110", "1010001101111110", "1010001101111110", "1010001101111110", "1010001101111101", "1010001101111111", "1010001001111111", "1010001001111111", "1010001001111111", "1010001101111111", "1010001101111111", "1010001101111111", "1010000101111110", "1001110001111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010001001111100", "1010001001111101", "1010000101111100", "1010001001111100", "1010001001111100", "1010001001111100", "1010001101111100", "1010010001111100", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010001101111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010001101111011", "1010001001111100", "1010001001111100", "1010001101111011", "1010001001111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010001001111100", "1010001101111100", "1010001001111100", "1010001101111100", "1010001001111100", "1010001101111100", "1010010001111011", "1010001101111100", "1010010001111011", "1010000101111100", "1010000101111101", "1010000101111100", "1010000001111101", "1010000101111101", "1010000101111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111101111101", "1010001001111101", "1010001001111101", "1010010001111101", "1010010001111110", "1010010001111110", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111110", "1010010101111101", "1010010101111101", "1010010101111110", "1010010101111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010001001111110", "1010001101111101", "1010001101111101", "1010000101111111", "1001110110000100", "1001100110000110", "1001011110000111", "1001101010000101", "1010000101111111", "1001111101111111", "1001111001111110", "1001111101111101", "1001111101111101", "1001111101111101", "1001111001111110", "1001110101111110", "1001110101111101", "1001110101111101", "1001111001111110", "1001111101111101", "1001111101111101", "1001111001111101", "1001010101111110", "1000011101111110", "0111111101111111", "0111111101111111", "0111111101111111", "1000000101111111", "1010001101111110", "1010001101111101", "1010001101111101", "1010001101111110", "1010001101111111", "1010001101111110", "1010001101111101", "1010001001111111", "1010001001111111", "1010001001111111", "1010001001111111", "1010001101111111", "1010001001111111", "1010001101111111", "1010010001111110", "1010001001111101", "1001110001111101", "1001100101111101", "1001100101111100", "1001101101111101", "1001101101111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000101111101", "1010000101111100", "1010000101111101", "1010001001111100", "1010001001111100", "1010001101111011", "1010001101111100", "1010001001111011", "1010001101111100", "1010001101111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111100", "1010010001111011", "1010010001111100", "1010010001111011", "1010001101111011", "1010000101111101", "1010000101111101", "1010000101111101", "1010001001111100", "1010001001111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010001001111100", "1010000101111100", "1010001101111100", "1010001001111100", "1010001001111100", "1010001101111011", "1010001001111100", "1010010001111011", "1010001001111100", "1010001001111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000001111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1010000101111101", "1010001001111101", "1010001101111101", "1010001101111101", "1010001101111110", "1010010001111110", "1010010001111101", "1010010001111110", "1010010001111111", "1010010001111110", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111110", "1010000010000001", "1001101010000110", "1001011110000110", "1001011110000111", "1001111010000100", "1010000001111111", "1001111101111111", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001110101111110", "1001110101111110", "1001110101111110", "1001110101111110", "1001111101111101", "1001111001111101", "1001010101111110", "1000011001111111", "0111111101111111", "0111111101111111", "1000000001111111", "1000000101111111", "1000001001111110", "1010001101111110", "1010001101111110", "1010001101111110", "1010001101111110", "1010001101111111", "1010001101111110", "1010001001111111", "1010001001111111", "1010001101111111", "1010001001111111", "1010001101111111", "1010001001111111", "1010001101111110", "1010010001111110", "1010001101111111", "1010001001111101", "1001110001111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000101111101", "1010000101111101", "1010000101111100", "1010001001111100", "1010000101111100", "1010000101111100", "1010001001111100", "1010000101111101", "1010001101111011", "1010001101111100", "1010010001111011", "1010001101111100", "1010001101111100", "1010001101111011", "1010001101111011", "1010010001111011", "1010001101111011", "1010010001111011", "1010001101111011", "1010000101111100", "1010000101111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010001001111100", "1010001001111100", "1010000101111100", "1010000101111101", "1010001101111100", "1010001001111011", "1010001001111100", "1010001101111011", "1010000101111100", "1010000101111101", "1010000101111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000001111101", "1010000101111101", "1001111101111101", "1001111101111101", "1001111101111100", "1001110101111101", "1001110001111101", "1001110001111101", "1001111101111101", "1010000101111101", "1010000101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010010001111110", "1010010001111110", "1010010001111110", "1010010001111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001001111111", "1001111010000100", "1001100010000110", "1001010110000111", "1001100010000111", "1001111110000001", "1010000001111110", "1001111001111110", "1001111001111110", "1001111101111101", "1001111001111110", "1001111001111110", "1001110001111110", "1001110101111110", "1001111001111101", "1001110001111101", "1001001101111110", "1000010101111110", "1000000001111111", "0111111101111111", "0111111101111111", "1000001001111110", "1000001001111110", "1000000101111111", "1010001101111101", "1010001001111111", "1010001001111111", "1010001101111111", "1010001101111111", "1010001101111110", "1010001001111111", "1010001001111111", "1010001001111111", "1010001101111111", "1010001101111111", "1010001001111111", "1010001001111111", "1010010001111110", "1010001101111110", "1010001001111110", "1001110001111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111100", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000101111101", "1010000101111100", "1010000101111100", "1010000101111101", "1010000101111100", "1010000101111100", "1010000101111100", "1010001101111011", "1010001101111100", "1010010001111011", "1010010001111011", "1010001101111100", "1010001001111100", "1010001101111011", "1010001101111100", "1010001101111100", "1010001101111100", "1010001001111100", "1010000101111100", "1010000101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111100", "1010001001111100", "1010001001111100", "1010001001111100", "1010001101111011", "1010001001111100", "1010000101111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1001111101111101", "1010000001111101", "1001111101111101", "1001111101111100", "1001110101111101", "1001110001111101", "1001110101111101", "1001111101111101", "1010000001111101", "1010000101111101", "1010001001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010010001111101", "1010001101111110", "1010010001111110", "1010010001111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010010101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010000110000000", "1001110010000110", "1001011110000111", "1001011010000111", "1001101010000101", "1010000001111111", "1001111001111111", "1001111001111110", "1001111101111101", "1001110101111110", "1001110101111101", "1001110101111110", "1001110101111110", "1001110001111110", "1001001001111110", "1000010001111110", "0111111101111111", "0111111101111111", "1000000101111111", "1000001001111110", "1000001001111110", "1000000101111111", "1000000101111111", "1010001001111110", "1010001101111110", "1010001001111111", "1010001101111110", "1010001001111111", "1010001001111111", "1010001101111111", "1010010001111110", "1010010001111111", "1010010001111111", "1010010001111111", "1010001001111111", "1010001101111111", "1010001101111110", "1010001101111110", "1010001001111101", "1001110101111101", "1001100101111101", "1001100101111100", "1001101001111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001111101111100", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111100", "1010000101111100", "1010001001111100", "1010001001111011", "1010001101111100", "1010001101111011", "1010001001111100", "1010001101111011", "1010001001111100", "1010001101111011", "1010010001111011", "1010001101111100", "1010001001111100", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111101", "1010000101111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000101111100", "1010000101111100", "1010000101111101", "1010000101111101", "1010001001111100", "1010001101111011", "1010001101111011", "1010001101111100", "1010001001111011", "1010000101111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111100", "1001111101111101", "1001111101111100", "1001111001111100", "1001110101111101", "1001110101111101", "1001111101111101", "1010000101111101", "1010000101111101", "1010001001111101", "1010001001111101", "1010001001111110", "1010001101111101", "1010001101111110", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010001101111101", "1010001101111101", "1010001101111110", "1010001101111111", "1001111110000100", "1001100010000111", "1001011010000111", "1001011010001000", "1001111010000100", "1001111101111111", "1001111001111110", "1001110101111110", "1001110101111110", "1001110001111101", "1001110001111110", "1001101101111110", "1001000101111111", "1000001101111111", "0111111101111111", "0111111101111111", "1000000001111111", "1000001101111101", "1000001001111110", "1000000101111111", "1000000101111111", "0111111101111111", "1010001001111110", "1010001001111111", "1010001001111111", "1010001001111110", "1010001001111110", "1010001001111111", "1010001101111111", "1010010001111110", "1010010001111111", "1010010001111111", "1010001101111111", "1010001101111111", "1010001001111111", "1010001101111111", "1010001101111111", "1010001001111101", "1001110101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111100", "1001111001111100", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000101111100", "1010001001111100", "1010001001111100", "1010001001111100", "1010001001111100", "1010001101111011", "1010001101111011", "1010001101111011", "1010001101111011", "1010010001111011", "1010001101111100", "1010010001111011", "1010010001111011", "1010001001111100", "1010001001111100", "1010001101111011", "1010001001111100", "1010000101111100", "1010000101111100", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000101111100", "1010000101111101", "1010001001111100", "1010001001111100", "1010001001111100", "1010001001111011", "1010001101111011", "1010010001111011", "1010010001111011", "1010001001111100", "1010000101111100", "1010001001111100", "1010000101111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111100", "1001111101111101", "1001111001111101", "1001110101111101", "1001110101111100", "1001110101111101", "1001111101111101", "1010000001111101", "1010001001111101", "1010000101111110", "1010000101111110", "1010000101111101", "1010001001111101", "1010001101111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111110", "1010001001111111", "1001110010000110", "1001011110000111", "1001011010000111", "1001100110000111", "1010000010000001", "1001111001111111", "1001110101111110", "1001110001111101", "1001110001111101", "1001101101111110", "1001000101111111", "1000001101111111", "0111111101111111", "0111111101111111", "1000000101111110", "1000001101111110", "1000001001111110", "1000000101111111", "1000000001111111", "0111111101111111", "0111111101111111", "1010001001111110", "1010001101111110", "1010001001111110", "1010001001111110", "1010001101111110", "1010001101111110", "1010010001111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010001101111111", "1010001101111111", "1010001101111111", "1010010001111110", "1010010001111110", "1010001001111101", "1001110001111101", "1001100001111101", "1001100101111100", "1001101101111100", "1001101101111101", "1001110001111100", "1001110001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110101111100", "1001111001111100", "1001111101111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000101111100", "1010000101111100", "1010000101111100", "1010001001111011", "1010010001111011", "1010001101111011", "1010001101111100", "1010001101111011", "1010001101111011", "1010001101111011", "1010001101111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010001101111011", "1010001001111011", "1010000001111100", "1001110001111100", "1001101101111100", "1001100001111101", "1001010001111101", "1001000101111101", "1001001001111101", "1001001101111101", "1001010001111110", "1001011101111101", "1001110001111101", "1001111101111101", "1010000101111100", "1010000101111101", "1010001001111100", "1010001001111100", "1010001001111100", "1010001101111011", "1010001101111100", "1010001001111100", "1010001001111011", "1010000101111100", "1010000101111101", "1010000101111100", "1010000101111101", "1010000101111100", "1010000001111101", "1001111101111101", "1001111101111100", "1001111001111100", "1001110101111100", "1001110101111100", "1001111101111101", "1010000001111101", "1010001001111101", "1010000101111111", "1010000101111110", "1010000101111101", "1010001001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010001101111101", "1010001101111101", "1010001101111110", "1010000110000010", "1001100110000110", "1001011010000111", "1001011010000111", "1001110110000100", "1010000001111111", "1001110101111111", "1001110001111110", "1001101101111101", "1001000001111111", "1000001101111111", "1000000001111111", "0111111101111111", "1000000101111111", "1000001001111110", "1000001001111110", "1000001001111110", "1000000101111111", "0111111101111111", "0111111101111111", "0111111101111111", "1010001001111110", "1010001001111111", "1010001001111111", "1010001001111110", "1010001101111110", "1010001101111110", "1010010101111101", "1010010101111101", "1010010001111101", "1010010001111110", "1010010001111111", "1010001101111111", "1010001101111111", "1010010001111110", "1010010001111110", "1010001101111101", "1001110101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001111001111100", "1001111101111100", "1001111101111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111100", "1010000101111100", "1010001001111011", "1010001001111100", "1010001101111011", "1010010001111010", "1010010001111011", "1010010001111011", "1010010001111010", "1010001101111011", "1010010001111011", "1010001101111011", "1010010001111100", "1010010001111010", "1010010001111010", "1001111101111100", "1001100101111100", "1001011101111100", "1001010101111101", "1001010101111100", "1001010101111101", "1001001101111101", "1001001101111101", "1001000101111101", "1001000001111101", "1001000001111101", "1001000101111101", "1001000001111101", "1000111101111110", "1000111101111111", "1001001101111111", "1001101001111101", "1001111101111101", "1010000101111100", "1010000101111100", "1010001001111100", "1010001101111011", "1010001001111100", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111100", "1010000001111101", "1010000101111100", "1001111101111101", "1001111001111101", "1001110101111101", "1001110101111100", "1001110101111100", "1001111101111101", "1010000001111101", "1010000101111101", "1010000101111110", "1010000101111110", "1010000101111110", "1010000101111101", "1010001001111101", "1010001001111110", "1010001101111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001001111111", "1001111010000100", "1001011110000111", "1001011010000111", "1001011110000111", "1001111110000010", "1001111101111110", "1001110001111111", "1001000101111111", "1000010001111111", "1000000001111111", "1000000001111111", "1000000101111111", "1000001001111110", "1000001001111110", "1000000101111111", "1000000101111111", "0111111101111111", "0111111101111111", "1000000101111111", "0111111101111111", "1010001001111110", "1010001001111111", "1010001001111111", "1010001101111111", "1010001101111111", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010001101111111", "1010001101111111", "1010010001111111", "1010010001111111", "1010010001111101", "1010001101111101", "1001110001111101", "1001100001111101", "1001100001111101", "1001100101111101", "1001101101111100", "1001101101111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110101111100", "1001111001111101", "1001111101111101", "1010000001111101", "1010000101111100", "1010000101111101", "1010000101111100", "1010000101111100", "1010000101111100", "1010001101111011", "1010001101111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010010001111011", "1010001101111011", "1010010001111011", "1010001101111011", "1010000101111011", "1001111101111100", "1001100101111100", "1001011101111101", "1001011101111101", "1001011001111100", "1001011101111100", "1001011001111101", "1001010101111101", "1001010001111101", "1001010001111101", "1001001001111101", "1001000001111101", "1001000001111101", "1001000001111101", "1001000101111110", "1001000001111110", "1001000001111111", "1000111101111111", "1000111001111111", "1001000001111111", "1001100101111101", "1010000001111101", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111101", "1010000101111100", "1010000101111101", "1010000101111101", "1010000101111101", "1010000001111101", "1001111101111101", "1001111001111100", "1001110001111101", "1001110001111101", "1001110001111101", "1001111101111101", "1010000101111101", "1010000101111101", "1010000101111110", "1010001001111110", "1010001001111101", "1010000101111101", "1010001001111101", "1010001001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010001101111101", "1010010001111101", "1010001101111110", "1010001101111101", "1010001101111101", "1010001101111110", "1010000101111111", "1001101110000101", "1001011010000111", "1001010110000111", "1001100110000111", "1001111101111111", "1001010101111111", "1000010101111111", "1000000101111111", "1000000101111111", "1000000101111111", "1000001101111101", "1000001001111110", "1000001001111110", "1000000101111111", "0111111101111111", "0111111101111111", "1000000101111111", "1000000001111111", "1000000101111111", "1010000101111110", "1010001001111110", "1010001101111110", "1010001001111111", "1010001101111110", "1010010001111101", "1010001101111100", "1010001001111101", "1010010001111101", "1010010001111110", "1010010001111111", "1010010001111111", "1010010001111111", "1010010001111111", "1010010001111101", "1010001001111101", "1001110001111101", "1001011101111101", "1001011101111101", "1001011101111101", "1001100101111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110101111100", "1001111001111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111100", "1010001001111100", "1010001101111011", "1010010001111011", "1010010001111011", "1010010001111010", "1010000101111100", "1001111001111011", "1001100101111100", "1001100101111100", "1001101001111101", "1001100101111101", "1001100101111101", "1001100101111100", "1001100001111101", "1001100101111101", "1001011001111101", "1001011101111101", "1001011001111101", "1001010101111101", "1001010001111100", "1001001101111100", "1001001101111101", "1001001001111101", "1001000001111101", "1001000101111110", "1001000001111111", "1000111101111111", "1000111101111111", "1000111001111111", "1000110101111111", "1000111001111111", "1001000101111110", "1001110001111101", "1010000001111101", "1010000101111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000001111101", "1001111101111101", "1001111001111101", "1001111001111100", "1001110001111100", "1001110001111100", "1001110001111101", "1001111001111101", "1010000101111101", "1010001001111101", "1010001101111101", "1010001001111110", "1010001001111110", "1010000101111101", "1010000101111101", "1010001001111101", "1010001001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010001101111101", "1010001101111110", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111110", "1001111110000010", "1001100010000110", "1001010010000111", "1001010010000111", "1001110010000010", "1000100101111111", "1000001001111110", "1000000101111111", "1000000101111111", "1000001101111110", "1000001101111110", "1000001101111101", "1000000101111111", "0111111101111111", "0111111101111111", "1000000101111111", "1000000101111111", "1000001001111110", "1000010001111101", "1010001001111110", "1010001001111110", "1010001101111110", "1010001101111110", "1010010001111101", "1010000101111101", "1001111001111101", "1010000001111101", "1010010001111101", "1010010001111110", "1010010001111111", "1010010001111111", "1010010001111111", "1010001101111111", "1010001101111110", "1010001001111110", "1001110001111101", "1001011101111101", "1001011001111101", "1001011101111101", "1001100001111101", "1001100101111100", "1001101001111100", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111100", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000101111101", "1010000001111101", "1010000101111100", "1010000101111100", "1010001001111011", "1010001001111100", "1010001001111100", "1001111101111110", "1001110001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001101001111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001100001111101", "1001011101111101", "1001011101111101", "1001011001111101", "1001010101111100", "1001010001111101", "1001010001111101", "1001001001111101", "1001001001111110", "1001000001111110", "1000111101111111", "1001000001111111", "1000111101111111", "1000111101111111", "1000111101111111", "1000111001111111", "1000110101111111", "1000110001111111", "1000111001111111", "1001011101111110", "1001111101111101", "1001111101111101", "1010000001111101", "1001111101111101", "1010000001111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1010000101111101", "1010001001111101", "1010001101111101", "1010001101111101", "1010001001111110", "1010001001111101", "1010000101111101", "1010000101111101", "1010001001111101", "1010001001111101", "1010010001111101", "1010001101111101", "1010001001111110", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010001101111110", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111110", "1010001101111101", "1010001101111110", "1010010001111101", "1010001001111111", "1001110110000100", "1001011110000111", "1001101010000100", "1000111110000001", "1000010001111110", "1000000101111111", "1000000101111111", "1000010001111101", "1000010001111101", "1000001101111110", "1000000101111111", "0111111101111111", "0111111101111111", "1000000101111111", "1000000101111111", "1000000101111111", "1000010001111101", "1000010101111101", "1010001001111110", "1010001001111110", "1010001101111110", "1010010001111101", "1010001001111101", "1001111001111101", "1001101001111101", "1001111101111101", "1010010001111101", "1010010001111110", "1010010001111111", "1010010001111111", "1010010001111111", "1010010001111111", "1010010001111101", "1010001001111101", "1001110001111101", "1001011001111101", "1001011001111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001101001111100", "1001101001111101", "1001101101111101", "1001110001111101", "1001110101111101", "1001111001111100", "1001111101111100", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000101111100", "1010000101111100", "1010000101111101", "1001110101111110", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001101001111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001100001111101", "1001011101111101", "1001011101111101", "1001010101111101", "1001010001111101", "1001001001111101", "1001000101111110", "1001000101111110", "1001000001111111", "1000111101111111", "1000111101111111", "1000111101111111", "1000111101111111", "1000111101111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000110101111111", "1001000001111111", "1001110001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110101111100", "1001110001111101", "1001110001111100", "1001110001111101", "1001111101111101", "1010000101111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010001001111101", "1010001001111110", "1010000101111110", "1010000101111101", "1010000101111101", "1010001001111101", "1010001101111101", "1010010001111101", "1010001101111110", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010001101111110", "1010010001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010010001111101", "1010001101111101", "1010001101111110", "1010000101111111", "1001111010000001", "1001000110000000", "1000010001111111", "1000001101111110", "1000001001111110", "1000010001111101", "1000010001111101", "1000001101111110", "1000001001111110", "0111111101111111", "1000000101111111", "1000001001111110", "1000000101111111", "1000001001111110", "1000010101111101", "1000010101111101", "1000010001111101", "1010001001111110", "1010001101111110", "1010001101111110", "1010001101111101", "1001111101111101", "1001101001111101", "1001100101111101", "1001111101111101", "1010001101111101", "1010010001111110", "1010010001111111", "1010010001111111", "1010001101111111", "1010001101111111", "1010001101111110", "1010000101111110", "1001110001111101", "1001011001111101", "1001011001111101", "1001011101111101", "1001100001111101", "1001100101111101", "1001100101111101", "1001101101111100", "1001100101111101", "1001101101111101", "1001110001111101", "1001110101111100", "1001111001111100", "1001111001111100", "1001111101111101", "1001111101111101", "1010000001111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000101111100", "1010000101111101", "1010000101111101", "1010000101111101", "1001111001111110", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001101001111101", "1001101001111101", "1001101001111101", "1001101001111101", "1001100101111101", "1001100101111101", "1001100001111101", "1001011101111101", "1001011001111101", "1001010001111101", "1001001101111101", "1001000101111110", "1001000001111111", "1001000001111111", "1000111001111111", "1000111001111111", "1000110101111111", "1000111001111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000101101111111", "1000110101111111", "1001011101111110", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1010000101111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010001101111101", "1010001001111101", "1001111101111101", "1001111101111101", "1010000101111101", "1010001001111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010001101111101", "1010010001111101", "1010001101111101", "1010001101111110", "1010010001111101", "1010010001111101", "1010001101111101", "1010010001111101", "1010001101111101", "1010001101111101", "1010000101111110", "1001000101111111", "1000001101111111", "1000001001111110", "1000001001111110", "1000010001111101", "1000010001111101", "1000010001111101", "1000001101111101", "1000000101111111", "1000000101111111", "1000010001111101", "1000000101111111", "1000001101111110", "1000011001111101", "1000011001111111", "1000011001111101", "1000110001111110", "1010001001111110", "1010001101111110", "1010001101111110", "1010001001111101", "1001110001111101", "1001100101111100", "1001101001111100", "1001111101111101", "1010001101111101", "1010010001111110", "1010010001111111", "1010010001111111", "1010001101111111", "1010001101111111", "1010001101111110", "1010000101111110", "1001110001111110", "1001011001111101", "1001011101111101", "1001011101111101", "1001100101111101", "1001101001111100", "1001101001111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010000101111100", "1010000101111110", "1001111101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001101001111101", "1001101001111101", "1001101001111101", "1001101001111101", "1001100101111101", "1001100001111101", "1001011101111101", "1001010101111101", "1001001101111110", "1001000101111111", "1000111101111111", "1001000001111111", "1000111101111111", "1000111101111111", "1000110101111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000101101111111", "1000011101111111", "1000010001111111", "1000000101111111", "1000001001111111", "1001001101111111", "1001110101111101", "1001111001111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1010000101111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010001101111101", "1010000101111101", "1001111001111101", "1001110001111101", "1001110101111101", "1010000101111101", "1010001001111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010001101111101", "1010001101111101", "1010000101111110", "1001010101111110", "1000010001111110", "1000000101111110", "1000000101111111", "1000010001111101", "1000010101111101", "1000010001111101", "1000010001111101", "1000000101111111", "1000001001111110", "1000010001111101", "1000000101111111", "1000001101111110", "1000010101111101", "1000011001111111", "1000011001111110", "1000101101111110", "1001100101111111", "1010001001111110", "1010001101111101", "1010001001111101", "1001111001111101", "1001100101111101", "1001100001111100", "1001101001111100", "1001111101111101", "1010001101111101", "1010010001111110", "1010010001111111", "1010001101111111", "1010001101111111", "1010001001111111", "1010001101111110", "1010000101111101", "1001110001111101", "1001011101111101", "1001011001111101", "1001100001111101", "1001100101111101", "1001101001111101", "1001100101111101", "1001101101111100", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000101111101", "1010000101111101", "1010000101111101", "1010001001111100", "1010000001111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001111101111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001101001111101", "1001101101111101", "1001101001111101", "1001101001111101", "1001011101111101", "1001011001111101", "1001001101111110", "1001000101111111", "1001000101111111", "1000111101111111", "1000111101111111", "1000111101111111", "1000110001111111", "1000111001111111", "1000110101111111", "1000100101111111", "1000010001111111", "1000010010000000", "1000001101111111", "1000001101111111", "1000010010000000", "1000000101111111", "1000001110000000", "1001100101111110", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1010000101111101", "1010010001111101", "1010010101111101", "1010011001111100", "1010010001111101", "1010001101111101", "1010000101111101", "1001110101111101", "1001100101111101", "1001100101111101", "1001111001111101", "1010000101111101", "1010001101111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010001101111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010010001111110", "1010010001111101", "1010010001111101", "1010010001111101", "1010001001111101", "1001100101111110", "1000011001111111", "1000000101111111", "1000000101111111", "1000010001111101", "1000011101111100", "1000010101111101", "1000010001111101", "1000000101111110", "1000001001111110", "1000011001111101", "1000001001111110", "1000001001111110", "1000010101111101", "1000010101111111", "1000011001111111", "1000101101111111", "1001011001111110", "1001110001111111", "1010001101111101", "1010001101111101", "1010000001111101", "1001101001111101", "1001100101111100", "1001100101111100", "1001100101111101", "1001111101111101", "1010001001111110", "1010010001111110", "1010010001111110", "1010010001111110", "1010010001111111", "1010001101111111", "1010001001111110", "1010000101111101", "1001110001111101", "1001011101111101", "1001011001111101", "1001100001111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001101001111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000001111101", "1010000101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001100101111101", "1001100001111101", "1001010101111101", "1001001001111111", "1001000101111111", "1000111101111111", "1000111101111111", "1001000001111111", "1000110101111110", "1000100001111111", "1000010001111111", "1000011001111111", "1000010001111111", "1000010010000000", "1000010101111111", "1000010001111111", "1000011101111111", "1000010010000000", "1000000110000000", "1000011101111111", "1001101001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001111001111101", "1010000101111101", "1010010001111101", "1010010101111101", "1010011001111100", "1010010001111101", "1010001101111101", "1010000101111110", "1001110001111110", "1001010101111101", "1001010001111101", "1001101001111101", "1001111001111101", "1010000101111101", "1010001101111101", "1010001101111101", "1010010001111101", "1010001101111110", "1010001101111101", "1010001101111110", "1010010001111101", "1010010001111101", "1010001101111101", "1010010001111101", "1010001101111101", "1001111101111101", "1000101001111111", "1000000101111111", "1000000101111111", "1000001101111110", "1000011001111101", "1000010101111101", "1000010101111101", "1000001001111110", "1000000101111111", "1000010101111101", "1000001001111110", "1000001001111110", "1000010101111101", "1000011001111111", "1000011001111111", "1000110001111110", "1001010101111110", "1001101001111111", "1001101101111111", "1010001101111101", "1010000101111101", "1001110001111101", "1001011101111101", "1001100101111100", "1001100101111100", "1001100101111101", "1001111101111101", "1010001101111101", "1010010001111101", "1010010001111111", "1010001101111111", "1010001001111111", "1010001101111111", "1010001001111110", "1010000101111110", "1001110001111101", "1001011101111101", "1001011001111101", "1001100001111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010000001111101", "1010000101111101", "1001111001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001101001111101", "1001100101111101", "1001011001111101", "1001010001111111", "1001001101111110", "1001000101111110", "1001000101111101", "1000110001111111", "1000010101111111", "1000010001111111", "1000011001111111", "1000011001111111", "1000011001111111", "1000010001111111", "1000010101111111", "1000010101111111", "1000010101111111", "1000010001111111", "1000001101111111", "1000000101111111", "1000110001111111", "1001110001111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001111001111101", "1010000101111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010001101111101", "1010000101111101", "1001110001111110", "1001010001111110", "1000111101111111", "1001011001111110", "1001110001111101", "1010000001111101", "1010001001111101", "1010001101111101", "1010001001111110", "1010001101111101", "1010001101111101", "1010001101111110", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010000101111101", "1001000101111110", "1000001101111110", "1000001001111110", "1000001001111110", "1000011101111100", "1000011001111100", "1000011001111100", "1000001101111110", "1000000101111111", "1000010101111101", "1000010001111101", "1000001001111110", "1000011001111101", "1000011001111110", "1000010001111111", "1000110001111101", "1001010001111101", "1001100101111111", "1001101101111111", "1001100101111111", "1010001001111101", "1001111101111101", "1001100101111101", "1001100001111101", "1001100101111100", "1001100001111101", "1001100101111101", "1001111001111101", "1010001001111101", "1010010001111101", "1010001101111111", "1010001101111111", "1010001101111111", "1010001101111110", "1010001001111110", "1010000001111110", "1001110001111101", "1001011101111101", "1001011001111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111100", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000101111101", "1001111101111101", "1001111001111101", "1001111001111101", "1001110101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001100101111101", "1001010101111110", "1001011001111101", "1001010001111101", "1000111001111111", "1000011101111111", "1000100010000000", "1000100001111111", "1000011001111111", "1000010001111111", "1000011001111111", "1000100001111111", "1000011101111111", "1000010101111111", "1000001101111111", "1000001110000000", "1000001101111111", "1000010001111111", "1000000101111111", "1000001001111111", "1001001001111111", "1001101001111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001111001111101", "1010000101111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010001101111101", "1010001001111101", "1001110001111101", "1001010001111110", "1000100101111111", "1001000101111111", "1001100001111101", "1001110101111101", "1010000101111101", "1010001001111101", "1010001101111101", "1010001101111101", "1010001001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001001111110", "1001011101111110", "1000010001111110", "1000000101111110", "1000001001111110", "1000010101111101", "1000010101111101", "1000011001111100", "1000010001111101", "1000000101111111", "1000010101111110", "1000010101111101", "1000001101111110", "1000011101111100", "1000011001111110", "1000010001111110", "1000100101111101", "1001010001111110", "1001100001111110", "1001101001111111", "1001101001111111", "1001101001111111", "1010000101111101", "1001101101111101", "1001011101111101", "1001100001111101", "1001100101111100", "1001100001111100", "1001100101111100", "1001110101111101", "1010001001111101", "1010010001111110", "1010001101111111", "1010001001111111", "1010001101111111", "1010001001111110", "1010001101111101", "1010000001111110", "1001101101111101", "1001011101111101", "1001011001111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000101111101", "1010000001111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001110101111110", "1001110101111110", "1001110001111101", "1001110101111101", "1001110001111101", "1001110001111110", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001100001111101", "1001011101111101", "1001010001111101", "1000111101111111", "1000100101111111", "1000100101111111", "1000011101111111", "1000011101111111", "1000100001111111", "1000100101111111", "1000100101111111", "1000011001111111", "1000011101111111", "1000011101111111", "1000011101111111", "1000011101111111", "1000010101111111", "1000010001111111", "1000010001111111", "1000010001111111", "1000001001111111", "1000100101111111", "1001011101111110", "1001101001111110", "1001101101111101", "1001110001111101", "1001111001111101", "1010000101111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010010001111101", "1010001001111101", "1001110001111110", "1001001101111110", "1000100101111111", "1000101001111111", "1001010001111101", "1001101101111101", "1001111101111101", "1010001001111101", "1010001101111101", "1010001101111101", "1010001101111101", "1010001001111110", "1010001101111101", "1010001101111101", "1010001001111110", "1001110101111110", "1000100001111110", "1000000101111111", "1000001001111110", "1000010101111101", "1000011001111100", "1000010101111101", "1000010001111101", "1000001001111110", "1000010001111110", "1000011001111110", "1000001101111110", "1000010101111101", "1000011001111101", "1000010101111111", "1000100001111110", "1001010001111101", "1001011101111111", "1001100101111111", "1001101001111111", "1001101001111111", "1001110001111111", "1001110101111101", "1001100001111101", "1001100001111100", "1001100001111101", "1001100001111101", "1001100001111101", "1001100101111101", "1001110101111101", "1010001001111101", "1010001101111110", "1010001001111111", "1010001001111111", "1010001001111111", "1010001001111110", "1010001001111110", "1010000001111110", "1001110001111101", "1001011101111101", "1001011001111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010001001111101", "1001111001111101", "1001110101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001110101111110", "1001110101111101", "1001111001111101", "1001111001111101", "1001111001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001101101111101", "1001100101111101", "1001010001111110", "1000110101111111", "1000110001111111", "1000101101111111", "1000110001111111", "1000110001111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000011101111111", "1000011101111111", "1000010101111111", "1000010101111111", "1000010001111111", "1000010101111111", "1000010101111111", "1000010110000000", "1000010010000000", "1000010110000001", "1000010010000000", "1000010101111111", "1001100001111110", "1001101001111110", "1001101101111101", "1001111001111101", "1010000101111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010001101111101", "1010001101111101", "1010000101111101", "1001110001111101", "1001010001111110", "1000100101111111", "1000100001111111", "1000111001111111", "1001011101111101", "1001110001111101", "1010000101111101", "1010001001111101", "1010001101111101", "1010001001111110", "1010001101111101", "1010001101111101", "1010001101111101", "1010000001111110", "1000111101111110", "1000001001111101", "1000000101111110", "1000010001111101", "1000011101111101", "1000011001111101", "1000011001111100", "1000001101111110", "1000010001111101", "1000011101111100", "1000010001111101", "1000010101111101", "1000011001111110", "1000010001111111", "1000010101111110", "1001000101111101", "1001011101111110", "1001100101111111", "1001100101111111", "1001101001111111", "1001101101111111", "1001110001111111", "1001100101111101", "1001011101111101", "1001100001111100", "1001100001111100", "1001100001111101", "1001100101111100", "1001100101111101", "1001110001111101", "1010001001111101", "1010001101111101", "1010001001111111", "1010001001111111", "1010001101111110", "1010001101111110", "1010001001111110", "1010000001111110", "1001110001111101", "1001011101111101", "1001011001111101", "1001011101111101", "1001100101111100", "1001100101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000101111111", "1010000101111101", "1001111001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001110101111110", "1001110101111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001100101111101", "1001001101111111", "1001001001111111", "1000110101111111", "1000110001111111", "1000111001111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000101101111111", "1000011101111111", "1000011101111111", "1000100001111111", "1000010101111111", "1000011101111111", "1000010101111111", "1000010110000000", "1000010101111111", "1000010110000000", "1000010001111111", "1000010101111111", "1000010010000000", "1000001110000000", "1000001110000000", "1000110001111111", "1001100101111110", "1001110001111101", "1001110101111101", "1010000101111101", "1010001101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010001001111101", "1010000101111101", "1001110001111101", "1001010001111110", "1000101001111111", "1000011101111111", "1000100101111111", "1001000101111111", "1001100101111110", "1001111101111101", "1010000101111101", "1010001001111101", "1010000101111110", "1010000101111110", "1010001001111101", "1010000101111101", "1001011001111110", "1000010001111110", "1000000101111111", "1000010001111101", "1000011001111101", "1000011001111101", "1000011001111101", "1000010001111101", "1000001101111101", "1000011001111100", "1000010001111101", "1000010001111101", "1000011101111111", "1000010101111111", "1000010101111111", "1000111001111101", "1001011101111110", "1001100101111110", "1001100001111111", "1001101001111111", "1001101101111111", "1001110001111111", "1001110001111111", "1001100101111100", "1001100001111101", "1001100001111100", "1001100001111100", "1001100001111101", "1001100001111101", "1001100101111101", "1001110001111110", "1010000101111101", "1010001001111110", "1010001001111111", "1010001001111111", "1010001001111111", "1010001101111101", "1010001001111110", "1010000101111101", "1001110001111101", "1001011001111101", "1001010101111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101101111100", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111110", "1010000101111111", "1001111101111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110101111110", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001011101111110", "1001010001111111", "1000111101111111", "1001000101111111", "1001001001111111", "1000111001111111", "1000110101111111", "1000111101111111", "1000110001111111", "1000101101111111", "1000101001111111", "1000100101111111", "1000011001111111", "1000010101111111", "1000011101111111", "1000010101111111", "1000010101111111", "1000010101111111", "1000011001111111", "1000010001111111", "1000010001111111", "1000011001111111", "1000010001111111", "1000001110000000", "1000000110000000", "1000000010000000", "1001001001111111", "1001101001111110", "1001110101111101", "1010000101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010000101111101", "1001110001111110", "1001010001111110", "1000101101111111", "1000100001111111", "1000011101111111", "1000101101111111", "1001010001111110", "1001100101111111", "1001011101111111", "1001000101111111", "1001010101111111", "1001101101111110", "1001111001111101", "1001101101111110", "1000100001111111", "1000000101111111", "1000001001111110", "1000011001111101", "1000011001111110", "1000011001111100", "1000010101111101", "1000001101111110", "1000010101111101", "1000010101111101", "1000010001111101", "1000011101111110", "1000011001111111", "1000011001111111", "1000110101111110", "1001011101111101", "1001100101111110", "1001100001111110", "1001100101111111", "1001101101111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001011101111101", "1001011101111101", "1001011101111100", "1001011101111101", "1001011101111101", "1001100001111100", "1001100101111100", "1001110001111101", "1010000101111101", "1010001101111101", "1010001001111111", "1010001001111111", "1010001001111111", "1010001001111111", "1010001001111110", "1010000101111101", "1001110001111101", "1001011001111101", "1001011001111101", "1001011101111101", "1001100101111100", "1001100101111101", "1001101001111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111111", "1010000101111111", "1001111101111101", "1001111001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001100101111110", "1001001001111111", "1001000101111111", "1001010001111111", "1001000101111111", "1000111101111111", "1001000101111111", "1001000101111111", "1000111101111111", "1000110001111111", "1000101001111111", "1000100101111111", "1000101001111111", "1000100001111111", "1000011001111111", "1000011101111111", "1000011101111111", "1000011001111111", "1000011001111111", "1000011101111111", "1000011001111111", "1000010001111111", "1000010001111111", "1000010001111111", "1000010001111111", "1000001110000000", "1000000001111111", "1000011001111111", "1001100101111101", "1001110101111101", "1010000101111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010000101111101", "1001110001111110", "1001010001111110", "1000110001111111", "1000100101111111", "1000100010000000", "1000100001111111", "1000110101111111", "1000100110000000", "1000011001111111", "1000100101111111", "1000011101111111", "1000011001111111", "1000100101111111", "1000110001111111", "1000001101111110", "1000001001111110", "1000010001111101", "1000011001111101", "1000010101111101", "1000011001111101", "1000010001111101", "1000010001111101", "1000010101111101", "1000010001111101", "1000011001111110", "1000011101111111", "1000011101111111", "1000110001111111", "1001010101111101", "1001101001111101", "1001100101111110", "1001100101111111", "1001101001111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001011001111101", "1001011001111101", "1001011101111101", "1001011101111101", "1001100101111100", "1001100101111100", "1001100101111100", "1001110001111101", "1010000101111101", "1010001001111110", "1010001001111111", "1010001001111110", "1010001001111110", "1010001001111110", "1010001001111110", "1010000101111101", "1001101101111101", "1001010101111101", "1001010101111101", "1001011001111101", "1001100001111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001100101111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111110", "1001111110000010", "1010001101111111", "1001111101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001111101111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001100101111101", "1001100001111101", "1001010101111111", "1001010001111111", "1001001101111111", "1001001101111110", "1001001101111110", "1001001001111110", "1001000001111111", "1001000001111111", "1000111101111111", "1000110001111111", "1000110001111111", "1000101101111111", "1000101001111111", "1000101001111111", "1000101001111111", "1000100101111111", "1000011101111111", "1000011101111111", "1000011001111111", "1000011001111111", "1000011001111111", "1000011001111111", "1000010001111111", "1000010001111111", "1000010101111111", "1000010001111111", "1000001101111111", "0111111101111111", "1001000101111111", "1001110001111101", "1010000001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010010001111101", "1010000101111101", "1001110101111101", "1001011001111110", "1000110101111111", "1000101101111111", "1000100110000000", "1000011110000001", "1000010110000001", "1000101001111111", "1000100001111111", "1000001010000000", "1000000110000001", "1000000110000001", "1000001010000000", "1000001101111111", "1000001101111111", "1000010001111101", "1000011001111101", "1000011001111110", "1000010101111101", "1000010101111101", "1000001101111110", "1000010101111101", "1000010001111101", "1000011001111101", "1000011101111111", "1000010101111111", "1000100101111111", "1001010001111101", "1001100101111110", "1001100101111110", "1001100101111111", "1001101001111111", "1001101101111111", "1001110001111111", "1001101101111111", "1001110001111111", "1001101101111111", "1001011101111101", "1001011101111101", "1001011101111101", "1001100001111101", "1001100101111100", "1001100101111100", "1001100101111101", "1001110001111101", "1010000101111110", "1010001101111101", "1010001001111110", "1010000101111111", "1010000101111111", "1010001001111110", "1010001001111110", "1001111101111110", "1001101101111101", "1001010101111110", "1001010101111101", "1001011001111101", "1001100001111101", "1001101001111101", "1001101001111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001111101111111", "1001111110000100", "1010010001111110", "1001111101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001111001111101", "1001110101111101", "1001110001111101", "1001100101111101", "1001011101111110", "1001010101111111", "1001011101111110", "1001011101111101", "1001001101111110", "1001010001111111", "1001001001111111", "1001010001111111", "1001000101111111", "1000111001111111", "1000111101111111", "1000111001111111", "1000110101111111", "1000101001111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000100001111111", "1000100101111111", "1000011101111111", "1000011101111111", "1000100001111111", "1000100001111111", "1000011101111111", "1000010001111111", "1000010101111111", "1000010001111111", "1000001101111111", "1000010001111111", "1000000101111111", "1000001101111111", "1001100101111101", "1010000001111101", "1010010001111101", "1010010101111101", "1010010101111101", "1010010001111101", "1010001101111101", "1010000101111101", "1001110101111110", "1001011001111110", "1000111001111111", "1000101101111111", "1000011110000000", "1000011110000001", "1000110101111111", "1000010101111111", "1000010010000001", "1000010001111111", "1000010010000000", "1000011110000000", "1000010010000000", "1000010010000000", "1000001101111111", "1000010101111110", "1000011001111101", "1000011001111101", "1000010101111101", "1000010001111101", "1000010101111101", "1000010001111101", "1000010101111101", "1000011101111111", "1000011101111111", "1000011101111111", "1001000101111101", "1001100001111110", "1001100101111110", "1001100101111110", "1001101001111110", "1001110001111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001101101111111", "1001101101111111", "1001011101111101", "1001011101111101", "1001011101111101", "1001100101111100", "1001100101111101", "1001100101111101", "1001101001111101", "1001110101111101", "1010000101111101", "1010001101111101", "1010000101111111", "1010001001111110", "1010000101111111", "1010000101111111", "1010001001111110", "1010000001111111", "1001101101111101", "1001011001111101", "1001010101111101", "1001011101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111110", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111111", "1010000110000011", "1010001101111110", "1001111001111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111001111101", "1001111101111101", "1001110101111101", "1001110001111101", "1001101101111101", "1001011101111110", "1001011101111110", "1001100001111101", "1001010001111110", "1001010001111110", "1001010001111111", "1001010001111111", "1001010001111111", "1001000101111111", "1001000001111111", "1000111001111111", "1000111101111111", "1000111101111111", "1000111101111111", "1000111101111111", "1000111001111111", "1000101001111111", "1000100101111111", "1000101101111111", "1000101001111111", "1000110001111111", "1000100001111111", "1000100101111111", "1000011001111111", "1000010101111111", "1000011001111111", "1000011101111111", "1000010101111111", "1000010101111111", "1000010001111111", "1000010001111111", "1000000101111111", "1000101001111111", "1001111101111101", "1010010001111101", "1010010101111101", "1010010101111110", "1010010001111101", "1010010001111101", "1010000101111110", "1001110001111111", "1001010101111111", "1000111001111111", "1000011010000000", "1000100110000000", "1000110101111111", "1000010010000000", "1000010110000001", "1000010110000000", "1000011101111111", "1000100001111111", "1000011101111111", "1000010001111111", "1000010010000000", "1000010010000001", "1000011010000000", "1000011001111110", "1000011001111101", "1000010001111101", "1000010001111101", "1000010101111101", "1000010001111101", "1000011001111110", "1000011101111111", "1000011101111111", "1000110101111110", "1001011101111101", "1001100101111110", "1001101001111101", "1001100101111110", "1001110001111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001101101111111", "1001110001111111", "1001100101111100", "1001100101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001110001111101", "1001101101111101", "1001111001111101", "1010000101111110", "1010001101111101", "1010000101111111", "1010000101111111", "1010000101111111", "1010000101111111", "1010001001111110", "1010000101111111", "1001110001111110", "1001011001111101", "1001011101111101", "1001100001111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111001111110", "1001111101111101", "1001111101111110", "1001111110000001", "1010000110000001", "1010001101111101", "1001111101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001100101111101", "1001101001111101", "1001011101111101", "1001010001111101", "1001011101111101", "1001011001111110", "1001001101111111", "1001010001111111", "1001001001111111", "1001001001111111", "1001000101111111", "1001000101111111", "1001000001111111", "1001001001111110", "1001001001111111", "1000111001111111", "1000111101111111", "1000110101111111", "1000101101111111", "1000101101111111", "1000101101111111", "1000100101111111", "1000101001111111", "1000011101111111", "1000111001111111", "1000110001111110", "1000100001111111", "1000100001111111", "1000011101111111", "1000010101111111", "1000010101111111", "1000010101111111", "1000010001111111", "1000000101111111", "1000100001111111", "1010000101111101", "1010010101111110", "1010010101111110", "1010010001111101", "1010010001111101", "1010000001111110", "1001100101111111", "1000110010000000", "1000011110000001", "1000110001111111", "1000100101111111", "1000010010000000", "1000010110000000", "1000011101111111", "1000100001111111", "1000100001111111", "1000011101111111", "1000010001111111", "1000010010000000", "1000011001111111", "1000010010000001", "1000010101111111", "1000011001111110", "1000010101111101", "1000010101111101", "1000010101111101", "1000010101111101", "1000011001111110", "1000011101111111", "1000010101111111", "1000100101111111", "1001010001111101", "1001100101111110", "1001100101111101", "1001100101111110", "1001101101111110", "1001110001111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001100101111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001110001111100", "1001111101111101", "1010001001111101", "1010001001111110", "1010000101111111", "1010000101111111", "1010001001111110", "1010001001111110", "1010001001111110", "1010000101111110", "1001110001111110", "1001011101111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111110", "1001110010000011", "1010001010000000", "1010001101111101", "1001111101111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001101101111101", "1001110101111101", "1001100101111101", "1001100001111101", "1001100101111101", "1001011001111110", "1001011001111110", "1001010001111111", "1001001001111111", "1001001001111111", "1001010001111110", "1001001001111111", "1001000101111111", "1001010001111110", "1001001001111111", "1001000101111111", "1001000101111111", "1000111101111111", "1001000001111111", "1000111001111111", "1000110001111111", "1000101101111111", "1000011101111111", "1000100101111111", "1000110101111110", "1001000101111110", "1000110101111111", "1000100101111111", "1000011101111111", "1000011101111111", "1000011101111111", "1000011101111111", "1000100001111111", "1000011101111111", "1000010001111111", "1000001101111111", "1001001001111111", "1010010001111110", "1010011001111101", "1010010001111101", "1010000001111110", "1001001101111111", "1000100110000000", "1000101010000000", "1000110001111111", "1000011101111111", "1000010110000000", "1000011110000000", "1000011101111111", "1000100001111111", "1000100001111111", "1000100001111111", "1000010101111111", "1000010101111111", "1000010101111111", "1000011001111111", "1000010010000000", "1000010101111111", "1000011001111101", "1000010101111101", "1000010101111101", "1000010001111101", "1000010101111101", "1000011101111111", "1000011101111111", "1000011101111111", "1001000101111110", "1001100101111101", "1001100101111110", "1001100101111101", "1001101001111110", "1001110001111111", "1001101101111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001101101111111", "1001101101111111", "1001101101111111", "1001100101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110101111100", "1001111101111101", "1010001101111101", "1010001001111101", "1010000101111111", "1010000101111111", "1010001001111111", "1010001001111111", "1010001101111110", "1010000101111110", "1001110001111110", "1001011101111101", "1001011101111101", "1001100001111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111111", "1001110110000100", "1010010001111111", "1010001101111101", "1010000001111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001100101111101", "1001101001111101", "1001100101111101", "1001100101111101", "1001010101111110", "1001001001111110", "1001010101111101", "1001011001111110", "1001010001111110", "1001000001111111", "1001010101111110", "1001010101111110", "1001001101111111", "1001010001111110", "1001000101111111", "1001000101111111", "1001001001111111", "1001000101111110", "1001000101111111", "1000110101111111", "1000110101111111", "1000110101111110", "1000111101111110", "1000111101111111", "1000110101111111", "1000111001111111", "1000110001111111", "1000101101111110", "1000100101111111", "1000101101111110", "1000100101111111", "1000011101111110", "1000100101111101", "1000100001111110", "1000011101111110", "1000100001111110", "1010001101111110", "1010010001111111", "1001100101111111", "1000101101111111", "1000101010000000", "1000111010000000", "1000101001111111", "1000011010000000", "1000011110000000", "1000011101111111", "1000100001111111", "1000100001111111", "1000011001111111", "1000011101111111", "1000011101111111", "1000010101111111", "1000010001111111", "1000010001111111", "1000011110000000", "1000010010000000", "1000011001111111", "1000010101111110", "1000010001111101", "1000010101111101", "1000010001111101", "1000011001111110", "1000011101111111", "1000100001111111", "1000111101111110", "1001100001111101", "1001100101111110", "1001101001111101", "1001100101111110", "1001110001111110", "1001110001111111", "1001110001111111", "1001101101111111", "1001110001111111", "1001101101111111", "1001101101111111", "1001101001111111", "1001101101111111", "1001100101111101", "1001101001111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110101111101", "1010000001111101", "1010001001111101", "1010001101111101", "1010000101111111", "1010001001111111", "1010001001111111", "1010001001111110", "1010001001111110", "1010000101111110", "1001110001111110", "1001100001111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111111", "1001110110000100", "1010001101111111", "1010010001111101", "1010000101111101", "1001111001111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001011101111101", "1001011101111101", "1001011001111101", "1001010001111101", "1001010001111101", "1001010001111110", "1001011101111101", "1001011001111110", "1001010001111111", "1001010001111111", "1001001101111111", "1001010001111111", "1001010001111110", "1001000101111111", "1001000001111110", "1000111001111111", "1000111101111111", "1001001101111101", "1001000001111111", "1000111101111111", "1000111101111111", "1000111101111111", "1000101101111111", "1000101101111110", "1000101001111111", "1000101001111110", "1000110101111101", "1000101001111110", "1000101101111101", "1000100101111101", "1000101001111101", "1000100101111101", "1000011101111101", "1001001001111110", "1000111101111111", "1000101010000000", "1000110101111111", "1000101101111111", "1000011101111111", "1000011010000000", "1000011110000000", "1000011101111111", "1000100001111111", "1000011101111111", "1000011001111111", "1000011101111111", "1000100101111111", "1000100101111111", "1000010101111111", "1000010001111111", "1000010101111111", "1000011110000000", "1000010101111111", "1000011001111111", "1000010101111101", "1000010101111101", "1000010001111101", "1000011001111101", "1000011101111111", "1000011101111111", "1000101101111110", "1001010101111101", "1001100101111101", "1001100101111110", "1001100101111110", "1001101001111110", "1001110001111110", "1001110001111111", "1001110001111111", "1001110001111111", "1001101101111111", "1001101101111111", "1001101101111111", "1001101101111111", "1001101101111111", "1001101001111101", "1001101001111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001111101111101", "1010001101111101", "1010001101111110", "1010001001111110", "1010000101111111", "1010000101111111", "1010001001111111", "1010001001111111", "1010000101111110", "1001110001111110", "1001011101111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001110101111111", "1001111010000101", "1010001101111111", "1010010001111101", "1010001001111101", "1010000001111101", "1001111101111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001111001111101", "1001110101111101", "1001110101111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001100001111101", "1001100101111101", "1001011101111101", "1001010101111101", "1001010001111110", "1001010001111110", "1001100001111101", "1001011101111110", "1001010001111111", "1001010101111110", "1001011001111110", "1001010101111111", "1001001101111110", "1001010001111101", "1001010001111110", "1001000101111110", "1001000001111110", "1001000001111110", "1001000101111111", "1001000001111110", "1000111101111110", "1000110101111110", "1000110001111111", "1000110001111110", "1000110001111101", "1000111101111101", "1000111101111101", "1000110101111101", "1000110001111101", "1000110001111101", "1000110001111101", "1000110101111100", "1000110001111101", "1000101001111111", "1000110001111111", "1000111110000000", "1000101101111111", "1000100101111111", "1000011010000000", "1000100101111111", "1000100001111111", "1000011101111111", "1000100101111111", "1000100001111111", "1000011101111111", "1000011101111111", "1000100001111111", "1000111001111111", "1000100101111111", "1000011101111111", "1000011001111111", "1000011101111111", "1000011010000000", "1000011010000000", "1000010101111111", "1000010101111101", "1000010101111101", "1000010001111101", "1000011101111111", "1000011101111111", "1000011101111111", "1001000001111101", "1001100101111101", "1001101001111101", "1001100101111110", "1001100101111111", "1001101001111111", "1001101101111111", "1001110001111111", "1001101101111111", "1001101001111111", "1001101101111111", "1001101101111111", "1001101101111111", "1001101101111111", "1001101101111111", "1001100101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001111101111101", "1010001101111101", "1010001101111110", "1010000101111111", "1010000101111111", "1010000101111111", "1010000101111111", "1010001001111110", "1010000101111110", "1001110001111110", "1001011101111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001111101111101", "1001111101111110", "1001110010000001", "1001111110000100", "1010001110000000", "1010010001111101", "1010010001111101", "1010001101111101", "1001111101111101", "1001111001111101", "1001111001111101", "1001110001111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001110001111101", "1001100101111101", "1001110101111101", "1001110001111101", "1001101101111101", "1001100001111101", "1001110001111101", "1001101001111101", "1001011101111101", "1001001101111101", "1001011101111101", "1001100101111101", "1001010101111110", "1001010101111110", "1001100001111101", "1001010101111110", "1001010101111110", "1001010001111110", "1001010001111110", "1001001101111110", "1001010001111101", "1001010101111110", "1001010001111110", "1001000101111111", "1001000101111110", "1000111101111110", "1001000101111111", "1000111101111101", "1000110001111110", "1000111101111101", "1001000001111101", "1000111001111101", "1000111101111101", "1001000001111100", "1000110001111101", "1000111101111100", "1001000001111101", "1000111001111111", "1000110001111111", "1000111101111111", "1000110001111111", "1000100101111111", "1000011101111111", "1000011110000000", "1000100001111111", "1000100101111111", "1000011101111111", "1000011101111111", "1000100001111111", "1000011101111111", "1000011001111111", "1000011101111111", "1001000001111110", "1001010001111110", "1000111001111110", "1000110001111111", "1000100101111111", "1000100101111111", "1000010110000001", "1000010101111111", "1000010101111101", "1000010101111101", "1000010001111101", "1000011001111101", "1000011101111111", "1000010101111111", "1000101101111111", "1001011001111101", "1001101001111101", "1001101001111101", "1001100101111110", "1001100101111111", "1001101001111111", "1001101001111111", "1001101101111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101101111111", "1001101001111111", "1001101101111111", "1001101101111111", "1001100101111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001111101111101", "1010010001111101", "1010010001111110", "1010000101111111", "1010001001111111", "1010000101111111", "1010000101111111", "1010001001111110", "1010000101111110", "1001110001111110", "1001011101111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111110", "1001111001111110", "1001111101111110", "1001110010000001", "1001111110000100", "1010010001111111", "1010010001111111", "1010010001111110", "1010010001111101", "1010000101111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001101001111101", "1001110101111101", "1001111001111101", "1001110001111101", "1001100101111101", "1001101101111101", "1001100101111101", "1001100001111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001011101111101", "1001011101111101", "1001011101111101", "1001011001111101", "1001011101111101", "1001010101111101", "1001011001111101", "1001011001111101", "1001011101111101", "1001011001111101", "1001010101111110", "1001010101111101", "1001010001111110", "1001010001111101", "1001001001111110", "1000111101111101", "1001000001111101", "1001000001111101", "1001000101111100", "1001000101111100", "1000111101111100", "1000111001111100", "1001000101111100", "1001000101111100", "1001000101111110", "1000111001111111", "1000111001111111", "1000111001111111", "1000100101111111", "1000100110000000", "1000100110000000", "1000101101111111", "1000101001111111", "1000100101111111", "1000100001111111", "1000011101111111", "1000100001111111", "1000011101111111", "1000011101111111", "1000011101111111", "1000110001111111", "1001010101111110", "1001010001111101", "1001010001111101", "1001010001111101", "1000110101111111", "1000011101111111", "1000010101111111", "1000010001111111", "1000010101111101", "1000010001111101", "1000010101111101", "1000011101111111", "1000010101111111", "1000100001111110", "1001001101111101", "1001101001111101", "1001101101111101", "1001101001111101", "1001100101111110", "1001101001111111", "1001101101111111", "1001101101111110", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101101111111", "1001100101111100", "1001100101111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001110101111101", "1001111101111101", "1010010001111101", "1010001101111110", "1010000101111111", "1010000101111111", "1010000101111111", "1010000101111111", "1010001001111110", "1010000101111110", "1001110001111110", "1001011101111101", "1001100001111101", "1001100101111101", "1001101001111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110101111100", "1001110101111101", "1001111001111101", "1001111101111110", "1001110010000010", "1010000110000011", "1010010010000000", "1010010001111111", "1010010001111111", "1010010001111101", "1010001101111101", "1001111001111101", "1001110001111101", "1001111001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001101001111101", "1001111001111101", "1001111101111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001100101111101", "1001100101111101", "1001100001111101", "1001101001111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001100001111101", "1001011001111101", "1001011101111101", "1001011001111101", "1001011101111101", "1001011101111101", "1001011101111101", "1001011001111110", "1001010101111101", "1001011001111110", "1001010101111101", "1001010101111101", "1001010001111101", "1001010001111101", "1001001001111101", "1001000101111100", "1001001001111101", "1001000101111100", "1001000101111100", "1001000101111100", "1001000101111011", "1001000101111101", "1000111101111111", "1001000001111111", "1000111101111111", "1000110001111111", "1000100001111111", "1000100101111111", "1000101101111111", "1000101101111111", "1000101001111111", "1000100101111111", "1000100101111111", "1000011101111111", "1000011101111111", "1000011101111111", "1000011101111111", "1000010101111111", "1000011101111111", "1001010001111101", "1001010001111101", "1001011001111110", "1001100001111110", "1001010001111101", "1000101101111111", "1000010110000000", "1000010101111111", "1000010101111101", "1000010101111101", "1000010001111101", "1000011101111110", "1000011101111111", "1000010101111111", "1000111001111101", "1001011101111101", "1001101101111101", "1001101001111101", "1001100101111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001100101111100", "1001100101111101", "1001100101111100", "1001100101111101", "1001101001111101", "1001101101111101", "1001110001111101", "1010000101111101", "1010010001111101", "1010001101111110", "1010000101111111", "1010000101111111", "1010000101111111", "1010000101111111", "1010001001111110", "1010000101111110", "1001110001111101", "1001011101111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001110110000011", "1010001010000100", "1010001110000001", "1010010101111111", "1010010101111110", "1010010001111101", "1010010001111101", "1010000101111101", "1001111101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001101101111110", "1001110101111101", "1001111001111110", "1001110101111101", "1001110101111101", "1001110001111101", "1001101101111101", "1001101001111101", "1001100101111100", "1001101101111101", "1001100101111101", "1001100101111100", "1001100101111101", "1001100101111101", "1001100101111101", "1001011101111100", "1001001101111011", "1001011001111101", "1001011001111101", "1001011001111101", "1001011001111101", "1001011101111101", "1001010101111101", "1001011101111101", "1001011001111101", "1001010101111101", "1001010001111101", "1001010001111100", "1001010001111100", "1001010001111100", "1001001101111011", "1001010001111011", "1001001101111011", "1001010001111100", "1001001001111111", "1001000101111111", "1001001001111111", "1000111001111111", "1000110010000000", "1000110001111111", "1000110101111111", "1000110001111111", "1000101101111111", "1000101001111111", "1000100101111111", "1000100001111111", "1000011001111111", "1000011001111111", "1000011101111111", "1000011101111111", "1000010101111111", "1000010101111111", "1000111101111110", "1001010001111101", "1001011001111110", "1001011101111101", "1001011101111101", "1001000101111110", "1000100001111111", "1000010101111111", "1000010101111111", "1000010101111110", "1000010101111101", "1000011001111101", "1000011101111111", "1000010001111111", "1000011101111110", "1001010001111101", "1001101001111101", "1001101101111101", "1001100101111110", "1001100101111111", "1001100101111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111101", "1001100101111101", "1001100101111101", "1001101001111100", "1001101001111101", "1001110001111101", "1001111001111101", "1010000101111101", "1010010001111101", "1010010001111110", "1010000101111111", "1010000101111111", "1010000001111111", "1010000101111111", "1010001001111110", "1010001001111110", "1001110101111110", "1001011101111101", "1001011101111101", "1001100101111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111001111110", "1001110010000100", "1010000010000101", "1010000110000011", "1010010010000000", "1010010101111111", "1010010101111110", "1010010101111101", "1010001001111101", "1001111001111101", "1010000001111101", "1001111101111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001110101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001100101111101", "1001100101111100", "1001011101111101", "1001001101111100", "1001000101111010", "1001000101111010", "1000111101111100", "1001000101111100", "1000111101111100", "1001010101111101", "1001011001111101", "1001011101111101", "1001010101111101", "1001010101111100", "1001011001111101", "1001010101111100", "1001011001111100", "1001010001111100", "1001010001111100", "1001010001111011", "1001010001111100", "1001010001111011", "1001010001111110", "1001000101111111", "1001001101111111", "1000111101111111", "1000110110000000", "1000110010000000", "1000110001111111", "1000110001111111", "1000101101111111", "1000101001111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000011101111111", "1000011001111111", "1000011001111111", "1000011001111111", "1000010101111111", "1000010001111111", "1000100001111111", "1001010001111101", "1001011101111101", "1001100001111101", "1001100101111101", "1001011101111110", "1000100101111111", "1000011101111111", "1000010001111111", "1000010101111111", "1000010101111111", "1000010101111101", "1000011001111111", "1000011101111111", "1000010001111111", "1000110101111101", "1001100101111101", "1001101001111101", "1001100101111110", "1001100101111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001101001111111", "1001101001111111", "1001101001111101", "1001101001111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001111101111101", "1010001101111100", "1010010001111101", "1010010001111110", "1010000101111111", "1010000101111111", "1010000101111111", "1010001001111111", "1010001101111110", "1010001001111110", "1001110101111101", "1001100001111101", "1001011101111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111001111101", "1001111101111110", "1001101110000100", "1001111110000110", "1010000010000011", "1010010010000000", "1010010001111111", "1010010001111111", "1010010101111111", "1010001101111101", "1010000001111101", "1001111101111101", "1001111001111101", "1001110101111101", "1001101101111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111001111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001101001111101", "1001101101111100", "1001011101111101", "1001010001111101", "1001011101111101", "1001011001111101", "1001001101111101", "1001000101111101", "1001000101111101", "1001010101111100", "1001000101111011", "1000110101111010", "1000111001111011", "1001000101111100", "1001010001111100", "1001000101111011", "1001000001111011", "1001000101111100", "1000111101111010", "1000110001111010", "1000101001111101", "1001010001111011", "1001011001111100", "1001010001111111", "1001010001111111", "1001001001111111", "1000101101111111", "1000110001111111", "1000110001111111", "1000101101111111", "1000101101111111", "1000101001111111", "1000101001111111", "1000100101111111", "1000100101111111", "1000100001111111", "1000011101111111", "1000011001111111", "1000011001111111", "1000010101111111", "1000011001111111", "1000010001111111", "1000011101111111", "1001001001111110", "1001011101111110", "1001100001111111", "1001101001111110", "1001100101111110", "1000111101111111", "1000100001111111", "1000010101111111", "1000010001111111", "1000010101111111", "1000010101111101", "1000010101111101", "1000011101111111", "1000010001111111", "1000011101111110", "1001010001111101", "1001100101111101", "1001101001111101", "1001100101111110", "1001100101111110", "1001100101111111", "1001100101111111", "1001101001111110", "1001101001111110", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001101001111101", "1001101101111100", "1001101001111101", "1001101001111101", "1001101101111101", "1001110101111100", "1010000001111101", "1010010001111100", "1010010101111101", "1010010001111110", "1010000101111111", "1010000101111111", "1010000101111111", "1010000101111111", "1010001001111111", "1010001001111110", "1001110101111110", "1001100001111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111100", "1001110101111101", "1001111101111101", "1001111101111110", "1001110010000100", "1001110110000110", "1001111110000100", "1010001110000010", "1010010001111111", "1010010001111111", "1010010001111111", "1010001001111110", "1001111001111101", "1001111001111101", "1001110101111101", "1001101101111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001100001111100", "1001011001111101", "1001011101111101", "1001010001111101", "1001001001111100", "1000111101111101", "1000100101111101", "1000011101111010", "1001001001111100", "1000101101111010", "1000100101111010", "1000010001111011", "1000000001111011", "1000000101111100", "1000010001111101", "1000100001111101", "1000100001111110", "1000001101111110", "1000010001111111", "1000010101111111", "1001000001111110", "1001010001111111", "1001011001111111", "1001000101111111", "1000110101111111", "1000110101111111", "1000110001111111", "1000101101111111", "1000101001111111", "1000101001111111", "1000101001111111", "1000100101111111", "1000100101111111", "1000100001111111", "1000011101111111", "1000011101111111", "1000010101111111", "1000011101111111", "1000011101111111", "1000011101111111", "1000110001111111", "1001010101111110", "1001100101111110", "1001100101111110", "1001101001111110", "1001101001111110", "1001010001111110", "1000101001111111", "1000011101111111", "1000010101111111", "1000010101111111", "1000010101111110", "1000010101111101", "1000011101111110", "1000011101111111", "1000010001111111", "1000110101111101", "1001100101111101", "1001100101111101", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001101001111110", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001101101111101", "1001101001111101", "1001101001111101", "1001101001111101", "1001101101111101", "1001110101111101", "1010000101111100", "1010010001111100", "1010010101111101", "1010010001111110", "1010000101111111", "1010000001111111", "1010000101111111", "1010001001111111", "1010001101111111", "1010001001111110", "1001110101111110", "1001100001111101", "1001011101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001110010000001", "1001111010000110", "1001111010000100", "1010000010000100", "1010010001111111", "1010010001111110", "1010001101111110", "1001111101111101", "1001111001111101", "1001110101111101", "1001101101111101", "1001110001111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001100101111101", "1001100101111101", "1001100101111100", "1001010001111100", "1001011001111101", "1001001101111101", "1001000001111100", "1000011101111100", "1000010001111100", "1000011101111011", "1000010001111010", "1000000101111101", "1000000101111110", "1000000101111101", "1000000001111101", "0111111101111101", "1000000001111110", "0111111101111111", "1000000101111111", "1000001001111111", "1000111101111111", "1001010001111111", "1001010101111111", "1000110101111111", "1000101101111111", "1000110001111111", "1000101101111111", "1000101101111111", "1000101101111111", "1000101001111111", "1000101101111111", "1000101001111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000011101111111", "1000011101111111", "1000100001111111", "1000100101111111", "1000111101111111", "1001011101111110", "1001100101111111", "1001101001111110", "1001100101111110", "1001101101111110", "1001101001111110", "1001011101111110", "1001001001111111", "1000100101111111", "1000011001111111", "1000010001111111", "1000011001111110", "1000010101111101", "1000010101111101", "1000011101111111", "1000010101111111", "1000010101111111", "1001010001111101", "1001100101111101", "1001100101111101", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001101001111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110101111101", "1010000001111101", "1010010001111100", "1010010101111110", "1010010001111110", "1010000101111111", "1010000101111111", "1010000101111111", "1010001001111111", "1010001101111111", "1010001001111110", "1001110101111110", "1001100001111101", "1001011101111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111110", "1001111101111101", "1001110110000000", "1001110010000111", "1001111010000110", "1001111110000100", "1010011001111111", "1010010101111101", "1010000101111110", "1001111101111110", "1001111101111101", "1001110001111101", "1001110001111101", "1001111101111101", "1001111101111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001101001111101", "1001100001111101", "1001101001111101", "1001010001111101", "1000111101111100", "1000110001111101", "1000100001111101", "1000010001111110", "1000010101111111", "1000010101111110", "1000000101111100", "1000000001111100", "1000010001111101", "1000010001111100", "1000010001111101", "1000000001111110", "0111111101111101", "1000000001111110", "1000000101111111", "1000001101111111", "1001000001111111", "1001011001111111", "1001001101111111", "1001000001111111", "1001000101111111", "1000110001111111", "1000101101111111", "1000110001111111", "1000110001111111", "1000101101111111", "1000101101111111", "1000101101111111", "1000101001111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000101101111110", "1001011101111101", "1001101001111110", "1001101001111111", "1001101001111110", "1001101101111110", "1001101101111101", "1001101101111110", "1001011101111111", "1001000001111111", "1000100101111111", "1000011001111111", "1000010101111111", "1000010101111110", "1000010101111101", "1000010101111101", "1000011001111111", "1000011101111111", "1000010001111111", "1000101101111110", "1001100001111101", "1001100101111101", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111100", "1001111101111101", "1010010001111100", "1010010101111101", "1010010001111111", "1010000101111111", "1010000101111111", "1010000101111111", "1010000101111111", "1010001001111111", "1010001001111110", "1001111001111101", "1001011101111101", "1001011101111101", "1001100101111100", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001111001111111", "1001110010000110", "1001111110000110", "1001111110000100", "1010010110000001", "1010010001111110", "1010000101111101", "1001111101111110", "1001111001111101", "1001110001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111100", "1001110101111101", "1001110101111101", "1001110001111101", "1001011101111101", "1001101001111101", "1001010101111101", "1000100101111110", "1000011001111110", "1000010001111101", "1000001101111110", "1000010001111111", "1000010101111111", "1000010101111100", "1000001001111100", "1000001101111101", "1000010001111110", "1000001001111101", "1000000101111101", "0111111101111101", "0111111101111101", "1000000001111111", "1000011001111111", "1001010001111111", "1001011101111111", "1001001101111111", "1001000101111111", "1001000101111111", "1000111101111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000101001111111", "1000101101111111", "1000101001111111", "1000100101111111", "1000100101111111", "1000101001111111", "1000110001111110", "1000110001111101", "1000110001111011", "1001010101111101", "1001110001111110", "1001110001111111", "1001110101111111", "1001111001111110", "1001110101111110", "1001101001111110", "1001001001111111", "1000100001111111", "1000011001111111", "1000010101111111", "1000010101111110", "1000010101111110", "1000010101111101", "1000010101111101", "1000011101111111", "1000010101111111", "1000010101111111", "1001001001111101", "1001100101111101", "1001100101111101", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111111", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1010000001111100", "1010010001111100", "1010010001111101", "1010001101111111", "1010000101111111", "1010000101111111", "1010000101111111", "1010000101111111", "1010001101111110", "1010001001111110", "1001110101111110", "1001100001111101", "1001011101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111001111101", "1001111101111110", "1001101010000100", "1001111110000110", "1001111110000100", "1010001010000011", "1010000101111111", "1010000101111101", "1001111101111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001100001111100", "1001100101111100", "1001110001111101", "1001110001111101", "1001011001111101", "1001000101111101", "1000011001111111", "1000011001111111", "1000001001111110", "1000000001111111", "1000000101111110", "1000001101111110", "1000010001111101", "1000100001111101", "1000010001111110", "1000010101111101", "1000001001111100", "1000000001111110", "0111111101111110", "1000000101111111", "0111111101111101", "1000100001111110", "1001011001111111", "1001011101111111", "1001000001111111", "1000111001111111", "1000111101111111", "1000111101111111", "1000111001111111", "1000111101111111", "1000111101111110", "1000111001111111", "1000111001111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000101001111111", "1000101001111111", "1000110001111111", "1000110101111110", "1000110001111100", "1000110001111011", "1000110001111010", "1001010001111011", "1001111001111110", "1010000001111111", "1010000001111111", "1001111101111111", "1001110001111111", "1001001101111111", "1000011101111111", "1000011001111111", "1000011001111111", "1000010101111110", "1000010101111101", "1000010101111110", "1000010101111101", "1000011001111110", "1000011101111111", "1000010001111111", "1000101001111101", "1001011101111101", "1001100001111110", "1001100101111101", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111110", "1001100001111111", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111111", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111101111101", "1010001101111100", "1010010101111101", "1010010001111111", "1010000101111111", "1010000001111111", "1010000001111111", "1010000101111111", "1010001101111111", "1010001001111110", "1001110101111110", "1001011101111101", "1001011101111101", "1001100101111100", "1001101001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001110010000001", "1001110010000111", "1001111110000110", "1010000110000010", "1001111101111111", "1010000101111111", "1001111101111101", "1010000001111101", "1001111101111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001100101111100", "1001001101111101", "1001001101111101", "1000111101111110", "1000011001111111", "1000011001111110", "1000010001111110", "1000001101111110", "1000001001111111", "0111111101111111", "1000001001111110", "1000010001111101", "1000010001111111", "1000010101111110", "1000010001111101", "1000000101111101", "0111111101111101", "0111111101111100", "0111111101111110", "1000100001111101", "1001011001111111", "1001100001111110", "1000111101111111", "1000111001111111", "1000110101111111", "1000111101111111", "1000111001111111", "1000111001111111", "1000111101111110", "1000111101111111", "1000111101111111", "1000110101111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000110101111110", "1001000001111110", "1000111101111110", "1000111001111101", "1000110001111100", "1000110001111010", "1000110101111010", "1001000101111010", "1001110001111101", "1001111101111110", "1001111101111111", "1001101101111111", "1001001101111111", "1000011101111111", "1000011001111101", "1000011001111111", "1000011001111101", "1000010101111101", "1000011001111101", "1000010101111101", "1000010101111101", "1000011101111111", "1000011001111111", "1000010101111111", "1001000101111101", "1001011101111110", "1001011101111101", "1001100101111110", "1001100101111110", "1001100001111111", "1001100101111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111110", "1001100101111111", "1001100101111111", "1001100101111110", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1010000101111100", "1010010001111101", "1010010001111111", "1010000101111111", "1010000010000000", "1010000001111111", "1010000101111111", "1010001001111111", "1010001001111110", "1001111001111110", "1001011101111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111110", "1001111101111111", "1001101010000100", "1001110010000111", "1001111010000010", "1001111110000000", "1001111101111111", "1010000001111101", "1001111101111101", "1001111101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001101101111101", "1001110001111100", "1001110101111101", "1001101101111100", "1001011101111101", "1000111101111110", "1000101001111111", "1000011101111111", "1000010101111111", "1000001001111101", "1000000101111111", "1000001101111101", "1000000001111111", "0111111101111111", "1000001101111111", "1000000101111111", "1000001001111110", "1000010101111110", "1000010001111101", "1000000101111101", "1000000101111101", "0111110101111010", "1000011101111101", "1000111101111101", "1001001101111111", "1001000001111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000110001111111", "1000111001111110", "1000111001111111", "1001000001111110", "1000111101111110", "1000111101111110", "1000110101111111", "1000101101111111", "1000110101111110", "1000111101111100", "1001010001111011", "1001100001111101", "1001001001111101", "1000111101111100", "1000110101111100", "1000110001111011", "1000111001111010", "1000111101111010", "1001100101111100", "1001111001111110", "1001101001111111", "1001000001111111", "1000010001111110", "1000010001111101", "1000011001111101", "1000011001111110", "1000011001111101", "1000011001111110", "1000011001111101", "1000010001111101", "1000011001111101", "1000011101111111", "1000010001111111", "1000100101111110", "1001010001111101", "1001010101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111110", "1001100101111111", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1010000001111101", "1010010001111101", "1010010001111110", "1010000101111111", "1010000001111111", "1010000001111111", "1010000101111111", "1010001101111111", "1010001001111110", "1001111001111110", "1001100001111101", "1001011101111101", "1001100001111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111110", "1001111101111111", "1001101010000110", "1001111010000011", "1001111010000010", "1001111101111111", "1010000101111101", "1001111101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001101001111101", "1001100101111100", "1001100001111100", "1001011001111011", "1001011001111011", "1001011101111101", "1001001001111110", "1001000001111110", "1000101101111111", "1000011101111110", "1000010001111110", "1000000101111111", "1000000001111111", "1000001001111101", "0111111101111111", "1000000101111111", "1000001001111111", "1000001001111111", "1000010001111111", "1000010001111110", "1000010001111101", "1000001001111101", "1000000101111100", "1000011001111100", "1000100101111011", "1001000001111101", "1000110101111110", "1000111101111111", "1000110001111111", "1000110001111111", "1000111001111111", "1000110101111111", "1000111101111110", "1000111101111111", "1000111101111110", "1000110101111111", "1000110001111110", "1000110001111101", "1000111101111100", "1001000101111011", "1000111101111011", "1001000101111010", "1001100001111011", "1001011101111100", "1001000001111101", "1000111001111100", "1000110001111100", "1000111001111011", "1000111101111011", "1001010101111100", "1001100001111110", "1001000001111111", "1000010001111110", "1000001001111110", "1000010001111101", "1000011001111101", "1000011001111101", "1000011001111101", "1000010101111111", "1000010101111101", "1000010101111101", "1000011001111110", "1000011001111111", "1000010001111111", "1000110101111110", "1001010001111111", "1001010001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111110", "1001100101111110", "1001101001111101", "1001101001111110", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111111", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111101111101", "1010001001111110", "1010001101111110", "1010000101111111", "1010000001111111", "1010000101111111", "1010000101111111", "1010001001111111", "1010001001111110", "1001111101111110", "1001011101111101", "1001011101111101", "1001100001111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111110", "1010000001111110", "1001101110000100", "1001101010000101", "1001110110000011", "1010000101111111", "1010000001111101", "1001111101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1001110101111101", "1001100101111101", "1001100101111011", "1000111101111101", "1000011101111111", "1000011101111111", "1000100001111111", "1000011101111110", "1000010101111110", "1000000101111111", "1000001001111110", "1000001101111110", "1000001001111110", "1000000101111111", "0111111101111111", "0111111101111111", "0111111101111111", "1000000101111111", "1000000101111111", "1000010101111110", "1000011101111101", "1000001001111011", "1000011001111010", "1000111001111011", "1001000101111111", "1001000001111111", "1000111001111111", "1000111101111111", "1001000001111111", "1000111101111110", "1000111101111111", "1000111101111111", "1000111001111111", "1000111001111101", "1000111001111101", "1000111001111100", "1000111101111011", "1000111101111100", "1000111101111011", "1000111101111011", "1001011001111010", "1001101001111101", "1001001001111101", "1000101101111101", "1000110001111101", "1000110001111100", "1000111101111010", "1001010001111011", "1001100001111101", "1000100001111110", "1000000101111111", "1000000101111110", "1000010101111101", "1000011001111101", "1000011001111110", "1000010101111110", "1000011001111101", "1000010101111101", "1000010101111101", "1000011101111111", "1000010101111111", "1000011101111110", "1001001001111110", "1001010001111111", "1001010101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001101001111101", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001110001111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110101111101", "1010001001111101", "1010001101111101", "1010000101111111", "1001111101111111", "1010000001111111", "1010000001111111", "1010001001111111", "1010001001111110", "1001111101111110", "1001011101111101", "1001011101111101", "1001100101111101", "1001100101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111100", "1001110001111101", "1001110001111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111110", "1010000001111110", "1001110010000011", "1001100010000110", "1001110110000100", "1010000101111110", "1001111101111101", "1001111001111100", "1001110101111101", "1001110001111101", "1001110001111101", "1001111001111100", "1001111101111100", "1001110001111101", "1001011001111101", "1001010001111101", "1000110001111111", "1000010101111111", "1000001001111111", "1000001101111110", "1000010001111111", "1000010101111110", "1000010001111110", "1000001001111110", "1000000001111111", "1000000001111101", "1000000001111111", "0111111101111111", "0111111101111111", "0111111101111111", "0111111101111111", "1000010001111111", "1001000001111101", "1001001101111101", "1000011101111010", "1000110101111101", "1001001001111111", "1000111101111111", "1000110101111111", "1000111101111110", "1001000001111110", "1001000101111101", "1000111001111110", "1000111001111110", "1001000001111101", "1001000101111100", "1001000001111101", "1000111101111101", "1000110101111101", "1000111101111011", "1001000001111100", "1000111101111011", "1000111101111100", "1001010101111010", "1001101101111100", "1001010101111101", "1000101101111110", "1000110001111101", "1000101101111101", "1000111101111010", "1001001001111011", "1001010001111110", "1000011101111110", "1000001001111110", "1000010001111101", "1000011001111101", "1000011001111101", "1000010101111110", "1000011001111110", "1000011001111101", "1000010101111101", "1000011001111101", "1000011101111111", "1000010001111111", "1000110001111101", "1001010101111111", "1001010001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100101111110", "1001100101111111", "1001100101111110", "1001100101111110", "1001100101111110", "1001101001111101", "1001101001111101", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110101111101", "1010001001111110", "1010001001111110", "1010000101111111", "1010000001111111", "1010000001111111", "1010000101111111", "1010001001111111", "1010001001111111", "1001111101111110", "1001100001111101", "1001011101111101", "1001100101111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111101", "1001111101111110", "1001111101111110", "1010000101111101", "1001110010000010", "1001100110000111", "1001110110000001", "1010000101111101", "1001111101111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1000110101111110", "1000011101111111", "1000011101111110", "1000010001111110", "1000000001111111", "0111111101111111", "1000001101111111", "1000010001111101", "1000010001111111", "1000000001111111", "0111111101111111", "1000000001111101", "1000000101111100", "1000001001111110", "0111111101111111", "0111111101111111", "1000001101111111", "1001011101111111", "1001010001111110", "1001010001111110", "1000100101111011", "1000101101111101", "1001000001111111", "1000110001111111", "1000110001111111", "1001000001111110", "1001000101111101", "1000111101111110", "1000110001111110", "1001001001111101", "1001011001111011", "1001010001111011", "1001000101111100", "1000111101111100", "1000111001111100", "1000111001111100", "1000111001111101", "1000111001111101", "1000110101111101", "1001001001111011", "1001101101111011", "1001011101111101", "1000101101111111", "1000100101111111", "1000101101111110", "1000111001111011", "1001000101111011", "1000110101111111", "1000010101111110", "1000000101111111", "1000010001111101", "1000011001111101", "1000011001111110", "1000010101111111", "1000010101111110", "1000010101111101", "1000010001111101", "1000011101111111", "1000010101111111", "1000011001111111", "1001000101111101", "1001010101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100101111111", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001101001111101", "1001100101111110", "1001100101111110", "1001101001111110", "1001101001111110", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1010001001111101", "1010001101111101", "1010000101111111", "1010000001111111", "1010000001111111", "1010000101111111", "1010001001111111", "1010001001111110", "1001111101111110", "1001100001111101", "1001011101111101", "1001100101111101", "1001101001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001111001111110", "1001111101111101", "1010000001111101", "1010000101111101", "1010000101111101", "1010000001111111", "1001100110000111", "1001111101111111", "1010000101111101", "1001111101111101", "1001110101111101", "1001110101111101", "1001111101111101", "1001110001111101", "1001010001111101", "1001010001111101", "1001000101111110", "1000110001111110", "1000011101111110", "1000010001111110", "1000000001111111", "1000001001111111", "1000000001111111", "0111111101111111", "1000010001111110", "1000010001111101", "1000001101111101", "1000000101111110", "0111111101111111", "1000000101111101", "0111111101111111", "0111111101111111", "1000000101111111", "1001100001111111", "1001101001111110", "1001010101111110", "1001011001111110", "1000111001111011", "1000011101111010", "1000110001111101", "1000110001111111", "1000111001111111", "1000111101111110", "1001000001111110", "1000111101111101", "1001011101111100", "1001100001111010", "1001010101111011", "1001001001111100", "1000111101111100", "1000111001111101", "1000110101111101", "1000111001111100", "1000110101111101", "1000101101111101", "1000101101111101", "1000111101111100", "1001100101111010", "1001101001111101", "1000111001111101", "1000011101111111", "1000101001111111", "1000101101111101", "1001000001111010", "1000110001111101", "1000011101111111", "1000010101111101", "1000011001111101", "1000011001111101", "1000011001111101", "1000010001111111", "1000011001111110", "1000010001111101", "1000010101111101", "1000011101111111", "1000010001111111", "1000100101111110", "1001010001111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001100001111110", "1001100101111110", "1001100101111110", "1001100101111110", "1001100101111111", "1001101001111110", "1001101101111110", "1001110001111101", "1001110001111100", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001111001111101", "1010001001111101", "1010001001111110", "1010000101111111", "1001111101111111", "1010000101111111", "1010000001111111", "1010001101111111", "1010001001111110", "1001111101111110", "1001100001111101", "1001011101111101", "1001100101111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111110", "1001111101111101", "1010000001111101", "1010000101111110", "1010001001111101", "1010000101111101", "1001100110000100", "1010000001111111", "1010000101111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001111001111101", "1001110001111101", "1001011101111101", "1000111001111110", "1000011101111101", "1000010001111110", "1000010101111101", "1000000001111111", "1000000101111111", "1000001101111111", "1000000101111111", "1000000101111111", "0111111101111111", "1000001101111110", "1000001101111110", "1000001001111101", "1000001001111101", "1000000101111100", "0111111101111111", "1000000101111111", "1001010101111111", "1001101101111111", "1001010101111111", "1001010001111111", "1001001001111111", "1000110101111100", "1000111101111100", "1000111001111111", "1000101001111111", "1000111101111110", "1000111101111101", "1001001001111101", "1001100101111010", "1001100101111010", "1001011101111011", "1001010001111100", "1001000001111011", "1000111101111100", "1000111101111100", "1000111001111100", "1000110001111101", "1000110001111101", "1000101001111101", "1000100101111101", "1000111001111101", "1001011001111011", "1001101101111100", "1001000101111110", "1000011001111101", "1000100001111111", "1000101001111101", "1000111101111011", "1000111001111101", "1000011001111110", "1000010001111110", "1000011001111101", "1000011001111110", "1000010101111110", "1000010001111111", "1000010101111101", "1000010001111101", "1000011001111110", "1000011101111111", "1000010101111111", "1000111101111110", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111110", "1001011001111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111110", "1001011101111111", "1001100101111110", "1001100101111110", "1001101001111110", "1001100101111111", "1001101001111111", "1001110001111110", "1001110001111101", "1001110001111100", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001111001111101", "1010000101111110", "1010001001111111", "1010000101111111", "1001111101111111", "1010000001111111", "1010000101111111", "1010001001111111", "1010001001111110", "1001111101111110", "1001100101111101", "1001100001111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000101111101", "1010000101111101", "1010001101111101", "1010010001111100", "1010000101111111", "1001111110000001", "1010000101111101", "1010000001111101", "1010000001111101", "1001111001111101", "1001110101111101", "1001100001111101", "1000110101111110", "1000010101111101", "1000001101111111", "0111111101111111", "1000000101111111", "1000010001111110", "1000000101111111", "1000001001111110", "1000000101111111", "1000000101111111", "1000000101111111", "1000000001111111", "1000000101111110", "1000001101111101", "1000000101111110", "1000000101111101", "1000000101111110", "1001010001111111", "1001101001111111", "1001011001111110", "1001011101111111", "1001000101111111", "1000111101111111", "1000110001111100", "1000111001111100", "1000110001111111", "1000110101111110", "1001000101111101", "1001010001111100", "1001100101111011", "1001100101111010", "1001100001111010", "1001011101111010", "1001010001111011", "1001000101111011", "1000111101111100", "1000111101111100", "1000110001111101", "1000110001111101", "1000110001111101", "1000100101111101", "1000100101111101", "1000101001111101", "1001001101111011", "1001101101111100", "1001010101111101", "1000100001111101", "1000011101111101", "1000100101111111", "1001000001111011", "1001000001111101", "1000011001111110", "1000010101111101", "1000011101111101", "1000011001111110", "1000010101111110", "1000010101111111", "1000010101111101", "1000010101111101", "1000011101111111", "1000011001111111", "1000100001111111", "1001010001111110", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111110", "1001011001111111", "1001010101111111", "1001011001111111", "1001011101111111", "1001011101111110", "1001011101111111", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111111", "1001101001111111", "1001110001111111", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110101111101", "1010000101111101", "1010001001111110", "1010000001111111", "1001111101111111", "1010000001111111", "1010000001111111", "1010001001111111", "1010001001111110", "1001111101111110", "1001100101111101", "1001100001111101", "1001100101111101", "1001101101111101", "1001110001111100", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001111101111110", "1010000001111101", "1010000101111101", "1010000001111101", "1010000101111101", "1010001001111101", "1010000001111110", "1010000101111101", "1010000101111101", "1001110001111100", "1001011001111011", "1001010001111101", "1000101101111111", "1000010001111110", "1000000001111111", "1000000101111110", "1000000101111111", "0111111101111111", "1000001001111111", "1000000101111110", "1000001101111110", "1000000101111111", "0111111101111111", "1000000101111111", "1000000101111111", "1000000101111111", "1000001001111101", "1000000001111111", "1000000001111111", "1000110001111101", "1001101001111111", "1001011101111110", "1001100101111110", "1001011101111110", "1001000001111111", "1000110001111111", "1000110101111110", "1000110101111101", "1000110101111110", "1001001001111101", "1001011001111011", "1001100101111010", "1001100101111010", "1001100001111010", "1001100001111010", "1001011101111010", "1001011001111010", "1001001001111100", "1001000001111101", "1000111101111101", "1000111101111101", "1000110101111101", "1000110101111100", "1000110001111101", "1000101001111101", "1000101001111101", "1001000101111100", "1001101001111011", "1001011101111101", "1000100101111110", "1000010001111101", "1000100101111111", "1000111101111100", "1001000001111101", "1000100001111111", "1000010101111101", "1000011101111110", "1000011001111111", "1000010101111111", "1000010101111110", "1000010001111101", "1000011001111101", "1000011101111111", "1000010101111111", "1000111001111101", "1001011101111111", "1001100001111111", "1001011101111111", "1001100001111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001101101111111", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1010000101111101", "1010001001111110", "1010000001111111", "1010000001111111", "1010000101111111", "1010000001111111", "1010001001111111", "1010000101111111", "1001111101111110", "1001100101111101", "1001100001111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010001001111101", "1010001101111100", "1010001001111110", "1001111001111111", "1010000101111111", "1010000101111110", "1001100101111100", "1001011101111011", "1001110001111100", "1001001001111101", "1000010101111101", "1000000101111111", "0111111101111111", "1000000101111101", "1000000101111111", "1000001001111110", "1000010001111110", "1000001001111110", "1000000101111111", "1000000101111111", "0111111101111111", "1000000101111111", "0111111101111111", "1000001001111110", "1000001001111110", "1000001001111111", "1000101101111110", "1001100001111111", "1001010101111110", "1001100101111110", "1001011101111111", "1001011001111101", "1000111101111111", "1000110001111111", "1000110001111110", "1000111101111101", "1001000101111101", "1001011101111011", "1001011101111010", "1001011101111010", "1001011101111010", "1001011101111010", "1001011101111010", "1001011101111010", "1001011101111010", "1001010001111011", "1001001001111100", "1001000101111101", "1001000001111100", "1000111101111100", "1000111101111100", "1000111101111100", "1000110001111101", "1000101101111101", "1000111101111100", "1001100101111011", "1001011101111101", "1000100101111110", "1000010001111101", "1000100101111111", "1000111001111101", "1001000101111100", "1000100101111111", "1000011101111111", "1000011001111101", "1000010101111111", "1000010001111111", "1000010101111110", "1000010101111101", "1000011101111111", "1000011101111111", "1000011101111111", "1001001001111101", "1001100001111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111110", "1001100101111111", "1001100101111111", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111100", "1001110001111101", "1001110101111101", "1010000101111101", "1010001001111110", "1010000101111111", "1010000001111111", "1010000001111111", "1010000101111111", "1010001001111111", "1010001001111110", "1001111101111110", "1001100101111101", "1001100001111101", "1001100101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001111101111101", "1010000001111101", "1001111101111101", "1010000101111110", "1010001001111101", "1001111110000000", "1001110101111111", "1001000101111111", "1001001001111111", "1001100101111110", "1001101101111111", "1001110001111101", "1001011101111101", "1000011101111110", "1000000101111101", "0111111101111111", "1000001001111101", "0111111101111111", "1000000001111111", "1000000101111111", "1000000001111111", "0111111101111111", "0111111101111111", "0111111101111111", "1000001001111111", "1000000101111111", "1000000101111101", "1000010001111110", "1000001101111101", "1000011101111111", "1001100101111111", "1001100001111111", "1001011001111111", "1001010101111111", "1001001001111111", "1001010101111110", "1000111001111111", "1000101001111111", "1000110101111101", "1001001101111101", "1001011001111101", "1001010001111100", "1001001101111100", "1001010001111011", "1001011001111010", "1001011101111010", "1001011001111010", "1001011101111010", "1001100001111010", "1001011101111010", "1001010101111011", "1001001001111100", "1001001001111100", "1001000101111101", "1001000101111100", "1001000101111101", "1000111101111101", "1000111101111100", "1001010001111010", "1001010101111100", "1000111101111111", "1000011001111101", "1000001001111110", "1000011101111111", "1000110001111101", "1001001001111011", "1000100101111111", "1000011101111111", "1000011001111110", "1000010101111111", "1000010101111111", "1000010001111101", "1000010101111101", "1000011001111111", "1000011001111111", "1000110001111110", "1001011001111110", "1001011101111111", "1001100001111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100001111111", "1001100001111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1010000101111110", "1010001001111110", "1010000101111111", "1010000101111111", "1010000001111111", "1010000101111111", "1010001001111111", "1010001001111110", "1001111101111110", "1001100101111101", "1001011101111101", "1001100101111101", "1001101101111101", "1001110001111100", "1001110001111101", "1001110101111101", "1001110101111101", "1001110101111101", "1001111001111101", "1001111101111101", "1010000001111101", "1010000001111101", "1010000101111101", "1010001001111101", "1010000001111111", "1001101001111111", "1001000101111111", "1001000101111111", "1001100101111101", "1001101101111111", "1001010001111101", "1000110001111111", "1000010001111110", "1000000101111101", "1000000101111111", "1000000101111101", "0111111101111110", "0111111101111111", "1000001101111110", "0111111101111111", "1000000101111111", "1000000001111111", "0111111101111111", "0111111101111111", "1000001101111110", "1000000101111101", "1000010001111101", "1000010001111101", "1001011101111111", "1001100001111111", "1001011101111111", "1001011001111111", "1000111101111111", "1001001101111110", "1001001001111110", "1000101101111111", "1000111101111101", "1001100101111101", "1001101001111100", "1001100101111101", "1001100101111100", "1001011101111100", "1001010001111101", "1001001101111101", "1001010001111100", "1001011101111011", "1001100101111010", "1001100101111010", "1001100101111010", "1001011101111011", "1001010001111100", "1001010001111011", "1001010001111011", "1001010001111011", "1001010001111011", "1001010001111011", "1001001101111100", "1001000101111101", "1001001101111101", "1001001101111101", "1000101101111110", "1000010101111101", "1000011101111111", "1000101101111101", "1001001001111011", "1000101001111111", "1000011101111111", "1000011001111111", "1000010001111111", "1000010101111110", "1000010101111101", "1000011001111110", "1000011101111111", "1000011101111111", "1000111101111110", "1001011101111111", "1001011101111111", "1001100101111111", "1001110001111111", "1001110001111111", "1001101101111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001100101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1010000101111101", "1010001001111110", "1010000101111111", "1010000001111111", "1010000001111111", "1010000101111111", "1010000101111111", "1010001101111101", "1001111101111110", "1001100101111101", "1001100001111101", "1001100101111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001111101111101", "1010000001111110", "1010000101111101", "1010000101111101", "1010001001111110", "1001110010000000", "1001100101111111", "1001001101111110", "1001101001111101", "1001010001111110", "1000110001111111", "1000011001111110", "1000000101111101", "1000001101111101", "1000000101111100", "0111111101111111", "1000000101111101", "0111111101111111", "1000001101111110", "0111111101111111", "1000001001111111", "1000000101111111", "1000000001111111", "1000000101111111", "1000001001111110", "1000010001111110", "1000001001111111", "1001000001111110", "1001100101111111", "1001010001111111", "1001011101111111", "1000111101111111", "1000110101111111", "1001001101111101", "1000110001111111", "1001000001111110", "1001100101111101", "1001100001111100", "1001011101111101", "1001001001111101", "1001011101111101", "1001010001111101", "1001011001111101", "1001100101111101", "1001100101111101", "1001101101111100", "1001110001111010", "1001110001111010", "1001110001111001", "1001100001111010", "1001010001111101", "1001010001111011", "1001010001111010", "1001011101111010", "1001011101111100", "1001010101111101", "1001010001111101", "1001000101111110", "1001001101111101", "1001000101111110", "1000101101111111", "1000011001111101", "1000011101111110", "1000110001111101", "1001000101111011", "1000110001111110", "1000011101111111", "1000010101111111", "1000010001111111", "1000010101111101", "1000010101111101", "1000011101111111", "1000011001111111", "1000100101111111", "1001010001111110", "1001011101111111", "1001100001111111", "1001101001111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001110001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100001111111", "1001100001111111", "1001100001111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001101001111101", "1001110101111101", "1010000101111110", "1010001001111110", "1010000101111111", "1010000001111111", "1010000001111111", "1010000001111111", "1010000101111111", "1010001001111110", "1001111101111110", "1001100101111101", "1001100001111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001100101111101", "1001110001111111", "1010000101111110", "1010000001111101", "1010000101111101", "1001111101111110", "1001101101111110", "1001000101111110", "1000100001111111", "1000010001111110", "1000010001111110", "1000000101111101", "1000001101111101", "1000000101111101", "1000000101111101", "0111111101111111", "1000001001111110", "0111111101111111", "1000000101111111", "0111111101111111", "0111111101111111", "1000000101111101", "1000000001111111", "1000010001111101", "1000011001111101", "1000010001111101", "1000100101111111", "1001100101111111", "1001010001111111", "1001100001111111", "1001001101111111", "1000101101111111", "1000111101111110", "1000111101111110", "1001000001111111", "1001001101111110", "1000111001111111", "1000101101111111", "1000011101111111", "1000010101111110", "1000011001111111", "1000010101111110", "1000101001111111", "1001010001111101", "1001110001111100", "1001110101111100", "1001111101111010", "1001111101111010", "1001111001111010", "1001100101111010", "1001010001111011", "1001000101111011", "1001010001111010", "1001010101111100", "1000110101111110", "1000011101111111", "1000010001111111", "1000010101111110", "1000011001111110", "1000100001111111", "1000011001111111", "1000010001111101", "1000011101111101", "1000110001111110", "1001001001111011", "1000110101111101", "1000011101111111", "1000010101111111", "1000010001111111", "1000010001111101", "1000010101111110", "1000011101111111", "1000011101111111", "1000110001111111", "1001011101111111", "1001100101111111", "1001100101111110", "1001100101111111", "1001101101111111", "1001110001111111", "1001101101111111", "1001101101111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100001111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001101101111101", "1001101001111101", "1001101001111101", "1001101001111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001110001111101", "1010000101111110", "1010001001111110", "1010000101111111", "1010000001111111", "1010000001111111", "1010000001111111", "1010000101111111", "1010001001111110", "1001111101111101", "1001100001111101", "1001011101111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101001111111", "1001110010000001", "1010000101111111", "1010001001111110", "1010001001111110", "1001101101111101", "1001011101111101", "1000111001111110", "1000011101111110", "1000010001111101", "1000011001111011", "1000001101111101", "1000000101111110", "1000001001111110", "1000000101111101", "0111111101111101", "0111111101111111", "1000000001111111", "1000000101111111", "1000000101111110", "0111111101111111", "0111111101111111", "0111111101111111", "1000000101111101", "1000001001111110", "1000011101111111", "1000011001111110", "1001010101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1000111001111111", "1000101101111111", "1000111101111110", "1001000101111110", "1001000101111110", "1000100101111111", "1000010101111111", "1000010001111110", "1000001001111111", "1000011101111110", "1000101001111101", "1000111001111101", "1000100101111111", "1000111001111111", "1001100001111101", "1001110101111100", "1010000001111010", "1010000001111010", "1001111101111010", "1001100101111010", "1001000101111100", "1000111101111100", "1001000101111101", "1000011101111111", "1000010001111110", "1000011101111101", "1000111001111101", "1000010001111111", "1000001001111110", "1000011101111101", "1000001001111111", "1000010101111101", "1000011101111110", "1000101101111111", "1001001001111010", "1000110101111101", "1000011101111111", "1000011001111111", "1000010101111111", "1000010101111101", "1000011101111110", "1000011001111111", "1000011101111111", "1001000101111110", "1001100001111111", "1001100101111110", "1001100101111111", "1001100101111111", "1001100101111111", "1001101101111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101101111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111110", "1001100001111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001101101111101", "1001101101111101", "1001101001111101", "1001101001111100", "1001100101111101", "1001100101111100", "1001100101111100", "1001101101111101", "1010000101111110", "1010001001111110", "1010000101111111", "1010000001111111", "1010000001111111", "1010000001111111", "1010000101111111", "1010001001111110", "1001111101111110", "1001100101111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111110", "1001100101111110", "1001101001111111", "1001111101111111", "1010000101111111", "1010000001111111", "1001110001111101", "1001000101111110", "1000011101111111", "1000010001111110", "1000010001111110", "1000000101111111", "1000001101111101", "1000000101111111", "1000001001111101", "1000000101111101", "1000000001111110", "0111111101111111", "0111111101111111", "0111111101111111", "1000000101111110", "1000000001111111", "0111111101111111", "0111111101111111", "1000000001111111", "1000000001111111", "1000001001111111", "1000110001111110", "1001011001111111", "1001001001111111", "1001010101111111", "1001000001111111", "1000100101111111", "1000110001111111", "1001000101111110", "1001011001111101", "1001000101111101", "1000110001111111", "1001000001111110", "1000100101111111", "1000011101111110", "1000100101111111", "1000011101111101", "1000110001111101", "1001010001111100", "1001011101111101", "1001100101111101", "1001110001111100", "1001111001111100", "1001111101111010", "1001111101111010", "1001100101111010", "1000110101111101", "1001000101111100", "1001000101111110", "1000100101111111", "1000011001111111", "1000011101111111", "1001000001111101", "1000111101111111", "1000010001111110", "1000001001111110", "1000001101111110", "1000010101111101", "1000100001111101", "1000101001111111", "1001000101111011", "1000111101111101", "1000100001111111", "1000010101111111", "1000010101111110", "1000010101111101", "1000011101111110", "1000011001111111", "1000100001111111", "1001010001111110", "1001100101111110", "1001100101111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001101101111101", "1001101101111101", "1001101001111101", "1001100101111101", "1001100101111101", "1001100101111100", "1001100001111101", "1001101001111101", "1010000101111110", "1010001001111110", "1010000101111111", "1010000001111111", "1001111101111111", "1010000001111111", "1010000101111111", "1010001001111110", "1001111101111101", "1001101101111101", "1001101001111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001110001111101", "1001110101111101", "1001110001111110", "1001011101111110", "1001001101111111", "1001010101111111", "1001100101111111", "1001100010000011", "1001010010000100", "1001000101111111", "1000011101111111", "1000001001111111", "1000010101111110", "1000010001111110", "1000001001111101", "1000001001111101", "1000001101111110", "1000010001111101", "1000000001111100", "1000000101111101", "0111111101111101", "0111111101111111", "0111111101111111", "0111111101111111", "1000000101111111", "1000000001111111", "1000000101111111", "1000000001111111", "1000000101111111", "0111111101111111", "1000001001111111", "1001011101111110", "1001001001111110", "1001010101111110", "1001001001111111", "1000101101111111", "1000101101111111", "1001001001111101", "1001100101111101", "1001100101111100", "1001011101111101", "1001001101111101", "1001010001111101", "1001010101111100", "1000110101111101", "1000110001111101", "1000101101111101", "1000111101111110", "1001100101111010", "1001110101111010", "1001111001111100", "1001110101111100", "1001110101111011", "1001111101111010", "1001111101111010", "1001010001111011", "1000100101111101", "1001010001111011", "1001011101111101", "1000111101111101", "1000101101111110", "1000110001111101", "1001001001111101", "1001001101111101", "1000100101111111", "1000011101111101", "1000010001111101", "1000010101111101", "1000100101111110", "1000101001111111", "1001001001111011", "1000110101111110", "1000100101111111", "1000011001111111", "1000010101111101", "1000010101111101", "1000011101111111", "1000010101111111", "1000110001111111", "1001011101111110", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100001111111", "1001100001111111", "1001100001111111", "1001100001111111", "1001100001111111", "1001100101111111", "1001101101111111", "1001101110000001", "1001101101111101", "1001101101111101", "1001101001111101", "1001100101111101", "1001100101111100", "1001100101111100", "1001100001111101", "1001101001111101", "1010000001111110", "1010001001111111", "1010000101111111", "1010000001111111", "1001111101111111", "1001111101111111", "1010000101111111", "1010001001111110", "1001111101111110", "1001101101111101", "1001101101111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001100101111111", "1001000001111111", "1001010001111111", "1001011101111111", "1001101101111111", "1001100101111111", "1001001110000001", "1000100110000001", "1000010101111110", "1000010001111101", "1000010001111100", "1000001001111100", "0111111101111110", "0111111101111111", "1000000101111110", "1000000101111101", "1000000101111101", "0111111101111011", "1000000101111011", "0111111101111100", "1000001001111110", "0111111101111111", "0111111101111111", "0111111101111111", "1000000001111111", "1000000001111111", "1000000001111111", "1000000101111111", "1000000101111111", "1001000101111111", "1001011101111110", "1001010001111111", "1001010101111111", "1000110101111111", "1000100101111111", "1001010001111101", "1001101101111100", "1001101101111100", "1001101101111100", "1001101001111011", "1001100101111011", "1001011101111011", "1001011101111011", "1001011101111010", "1001011101111010", "1001010001111010", "1001010001111000", "1001001101110111", "1001100101111001", "1001111001111010", "1001110101111011", "1001111001111011", "1010000001111010", "1001111101111001", "1001001001111010", "1000010101111101", "1001001001111010", "1001010101111010", "1001011101111010", "1001011101111011", "1001010101111010", "1001010101111101", "1001000001111110", "1000110101111111", "1000101001111111", "1000011101111110", "1000011101111101", "1000101001111111", "1000101001111111", "1001001001111010", "1000111101111100", "1000100101111110", "1000011001111111", "1000010001111101", "1000011001111101", "1000011101111111", "1000011101111111", "1001000101111110", "1001100101111110", "1001100101111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111110", "1001100101111111", "1001101001111111", "1001101101111111", "1001110010000000", "1001110110000001", "1001110110000010", "1001110010000010", "1001110001111101", "1001110001111101", "1001101101111101", "1001100101111101", "1001100101111101", "1001100001111101", "1001011101111101", "1001101001111101", "1010000001111110", "1010001001111110", "1010000101111111", "1010000001111111", "1001111110000000", "1010000010000000", "1010000101111111", "1010001101111110", "1010000101111110", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001111101111110", "1001101001111111", "1001011101111111", "1001101101111111", "1001100101111111", "1001001101111101", "1001001001111110", "1000100101111111", "1000011001111110", "1000010001111111", "1000000001111011", "1000000101111101", "1000000101111100", "0111111101111110", "1000000101111111", "1000000101111110", "1000000001111101", "1000000001111110", "1000000001111011", "0111111101111010", "0111111101111011", "0111111101111110", "0111111101111111", "0111111101111111", "0111111101111111", "0111111101111111", "0111111101111111", "1000000101111111", "1000000101111111", "1000100001111110", "1001101001111111", "1001011001111111", "1001011101111111", "1001000001111111", "1000100101111111", "1001010001111101", "1001101101111100", "1001101101111011", "1001110001111011", "1001110001111010", "1001110001111010", "1001101101111011", "1001101001111011", "1001101101111011", "1001101001111011", "1001100101111010", "1001100001111010", "1001010101111010", "1001100001111001", "1001101001111001", "1001110001111010", "1001111001111010", "1001111101111010", "1010000101111001", "1001111101111001", "1001010101111001", "1000010101111100", "1001000101111001", "1001100001111001", "1001101001111010", "1001100101111011", "1001100001111011", "1001010001111101", "1001001101111101", "1001000101111101", "1000110101111111", "1000011101111110", "1000100101111110", "1000110001111111", "1000100101111111", "1001001101111011", "1000111101111100", "1000100101111111", "1000011001111111", "1000010101111101", "1000011101111110", "1000011101111111", "1000100101111111", "1001010101111111", "1001100101111110", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001101101111111", "1001110110000000", "1001111110000011", "1001111110000100", "1001111010000100", "1001111010000100", "1001110110000100", "1001101101111101", "1001101001111101", "1001100101111100", "1001100001111101", "1001011101111101", "1001011101111101", "1001011001111101", "1001100101111101", "1001111101111110", "1010001001111110", "1010000101111111", "1010000101111111", "1010000001111111", "1001111110000000", "1010000101111111", "1010001101111110", "1010000101111110", "1001101101111110", "1001101101111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001111001111111", "1001110001111111", "1001101001111101", "1001001101111101", "1000100101111111", "1000100101111110", "1000010101111110", "1000001001111110", "1000010001111110", "1000001001111101", "0111111101111011", "0111110101111010", "0111111101111101", "1000000101111111", "1000001101111110", "1000000101111101", "1000000001111011", "1000000001111101", "0111111101111100", "0111111101111100", "1000001001111110", "1000000101111111", "0111111101111111", "0111111101111111", "0111111101111111", "0111111101111111", "1000000101111111", "1000001101111110", "1001011001111111", "1001100101111111", "1001011101111111", "1001001001111111", "1000100101111111", "1001000101111110", "1001101101111101", "1001110001111011", "1001110001111011", "1001110001111011", "1001110001111010", "1001101101111010", "1001101001111010", "1001101001111010", "1001101101111010", "1001101001111010", "1001100101111010", "1001100001111010", "1001100001111001", "1001100101111000", "1001101001111001", "1001110101111010", "1001111101111001", "1010000001111001", "1010000101111001", "1010000101110111", "1001011101111000", "1000011001111011", "1000110101111010", "1001010001111001", "1001100101111001", "1001101101111010", "1001101101111100", "1001101101111100", "1001011101111101", "1001010101111101", "1001000001111110", "1000100101111111", "1000101001111111", "1000110001111111", "1000100101111111", "1001010001111011", "1001000101111011", "1000100101111111", "1000011001111111", "1000011001111101", "1000011101111111", "1000011001111111", "1000110001111111", "1001011101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001110001111111", "1001111010000011", "1001111010000101", "1001111110000101", "1010000010000101", "1001111110000100", "1001111110000100", "1001111010000100", "1001100101111101", "1001100101111101", "1001100001111101", "1001011001111101", "1001011001111101", "1001011001111101", "1001010101111101", "1001100001111101", "1001111101111101", "1010001001111110", "1010000101111111", "1010000001111111", "1010000010000000", "1010000010000000", "1010000101111111", "1010001001111110", "1010000101111110", "1001110001111101", "1001101001111101", "1001110001111101", "1001110001111110", "1001111001111101", "1001111101111101", "1001110101111101", "1001011101111101", "1001011101111101", "1000100101111100", "1000010101111011", "1000010001111110", "1000010101111110", "1000010101111101", "1000001001111101", "1000000101111011", "1000000101111101", "1000001001111101", "0111111101111111", "1000000001111111", "1000000101111110", "1000001001111101", "1000000001111101", "0111111101111010", "1000000101111100", "0111111101111010", "1000001101111110", "1000010001111110", "1000000101111111", "0111111101111111", "0111111101111111", "1000000001111111", "1000000101111111", "1000110101111110", "1001100101111111", "1001011001111110", "1001010001111111", "1000110101111111", "1000110001111111", "1001100001111101", "1001110001111100", "1001110101111011", "1001111001111010", "1001111101111010", "1001111001111001", "1001110001111000", "1001100101111001", "1001100101111010", "1001100001111001", "1001100101111001", "1001100001111001", "1001100101111001", "1001100101111001", "1001101001111001", "1001110001111001", "1001111101111001", "1001111101111001", "1010000001111001", "1010000101111000", "1010000101111000", "1001011101110111", "1000011101111010", "1000110001111010", "1001001101111001", "1001100001111001", "1001110001111010", "1001110001111010", "1001101101111011", "1001100101111100", "1001011101111100", "1000111101111110", "1000100101111111", "1000101101111111", "1000110101111111", "1000100101111111", "1001001101111100", "1001001001111011", "1000100101111111", "1000011001111111", "1000011001111110", "1000011101111111", "1000011001111111", "1001000101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111111", "1001100101111111", "1001100101111111", "1001110010000000", "1001111010000100", "1001111110000110", "1010000110000111", "1010000110000110", "1010000110000110", "1010000010000100", "1001111110000100", "1001111010000100", "1001100001111101", "1001011101111101", "1001011101111101", "1001011001111101", "1001011001111101", "1001010101111101", "1001010001111101", "1001011101111101", "1001111101111101", "1010000101111110", "1010000101111111", "1010000001111111", "1001111110000000", "1010000010000000", "1010000101111111", "1010001101111110", "1010000101111110", "1001110001111101", "1001101101111101", "1001110001111101", "1001110001111110", "1001110001111101", "1001100001111100", "1001000101111010", "1001001001111010", "1000100101111101", "1000010001111101", "1000010001111111", "1000010001111111", "1000011001111111", "1000001101111101", "1000000101111101", "1000000001111100", "1000000101111011", "0111111101111110", "0111111101111111", "0111111101111111", "0111111101111111", "1000000101111111", "1000001001111101", "1000010001111100", "0111111101111101", "1000010001111110", "1001001101111110", "1000111101111111", "1000000101111111", "0111111101111111", "0111111101111111", "1000000101111111", "1000010001111110", "1001011101111111", "1001100001111111", "1001010001111111", "1000111101111111", "1000011101111111", "1001000101111110", "1001100001111101", "1001110001111100", "1001111001111011", "1001111101111010", "1001111101111001", "1001111101111001", "1001110101110111", "1001101101111000", "1001100101111001", "1001100101111001", "1001100101111010", "1001100101111001", "1001100101111001", "1001100101111010", "1001110001111000", "1001111001111000", "1001111101111001", "1001111101111001", "1010000001111001", "1010000001111001", "1010000101111001", "1001100101110111", "1000011001111010", "1000101101111010", "1001010001111010", "1001100001111010", "1001110001111010", "1001110101111010", "1001101101111011", "1001100101111010", "1001011101111011", "1001000001111110", "1000101001111111", "1000110001111111", "1000110101111111", "1000100101111111", "1001001101111100", "1001010001111010", "1000101001111111", "1000011001111110", "1000011101111111", "1000011101111111", "1000100001111111", "1001010101111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100001111111", "1001100101111111", "1001100001111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001110001111111", "1001111110000100", "1010000010000110", "1010000110000111", "1010000110000111", "1010000110000110", "1010000110000110", "1010000010000101", "1001110110000101", "1001101110000100", "1001011001111101", "1001010101111101", "1001010101111101", "1001010001111101", "1001010101111101", "1001010101111101", "1001010001111110", "1001011101111101", "1001111101111110", "1010000101111110", "1010000101111111", "1010000001111111", "1010000001111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000101111110", "1001101101111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110101111101", "1001011001111101", "1000110001111101", "1000100001111110", "1000011101111101", "1000011101111111", "1000010101111110", "1000001101111101", "1000000101111101", "1000000101111011", "0111111101111101", "0111111101111101", "0111111101111111", "0111111101111111", "0111111101111111", "0111111101111111", "0111111101111111", "1000010001111111", "1000011101111111", "1000010001111111", "1000100101111111", "1001010101111111", "1001000001111111", "1000010001111111", "0111111101111111", "0111111101111111", "0111111101111111", "1000111101111111", "1001100101111111", "1001010001111111", "1001001101111111", "1000100101111111", "1000100001111111", "1001001001111101", "1001100101111100", "1001110001111100", "1001111101111010", "1001111101111010", "1010000101111001", "1010000001111001", "1001111101111000", "1001110001111000", "1001101101111001", "1001100101111001", "1001100101111001", "1001100101111001", "1001101001111001", "1001101001111001", "1001110001111001", "1001110101111001", "1001111101111001", "1001111101111001", "1010000001111001", "1010000101111001", "1010000101111000", "1001101001110111", "1000011101111010", "1000100101111010", "1001010101111010", "1001100101111010", "1001110001111001", "1001110101111010", "1001110001111011", "1001100001111010", "1001011101111011", "1001000001111110", "1000100101111111", "1000110001111111", "1000111101111110", "1000100101111111", "1001001001111101", "1001010001111011", "1000110001111110", "1000011001111111", "1000100001111111", "1000011101111111", "1000110001111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100001111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001101101111111", "1001111110000011", "1010000110000110", "1010001010000111", "1010000110000111", "1010000110000111", "1010000110000110", "1010000010000110", "1001110110000110", "1001100110000101", "1001011010000101", "1001010101111101", "1001010001111101", "1001001101111110", "1001001101111110", "1001010001111110", "1001001101111110", "1001001101111111", "1001011101111101", "1001111101111110", "1010000101111110", "1010000001111111", "1001111101111111", "1001111101111111", "1010000001111111", "1010000101111111", "1010001001111110", "1010000001111110", "1001101101111101", "1001100101111101", "1001101101111101", "1001110101111101", "1001111001111101", "1001111001111101", "1001010001111101", "1000100101111010", "1000011101111101", "1000110101111101", "1000100001111110", "1000010001111101", "1000001001111101", "1000001001111101", "0111110101111011", "0111111101111101", "1000000001111111", "1000000001111111", "0111111101111111", "0111111101111111", "0111111101111111", "0111111101111111", "1000000001111111", "1000010001111111", "1000011101111111", "1000111001111110", "1001000101111110", "1001010101111111", "1000100101111111", "0111111101111111", "1000000101111111", "1000011001111111", "1001100001111111", "1001011101111111", "1001000101111111", "1000110001111111", "1000011001111111", "1000101001111110", "1001000101111110", "1001100101111100", "1001110001111100", "1001111101111010", "1001111101111010", "1010000101111010", "1010000101111010", "1010000001111000", "1001111101111000", "1001110001111000", "1001101101111001", "1001101001111001", "1001100101111001", "1001101001111001", "1001101101111001", "1001110101111001", "1001111101111010", "1001111101111010", "1010000001111001", "1010000001111001", "1010000101111000", "1010000101111000", "1001111001110111", "1000110001111001", "1000011001111011", "1001010101111010", "1001100101111001", "1001101101111010", "1001110001111010", "1001101101111010", "1001100101111010", "1001011101111100", "1000111001111110", "1000100101111110", "1000101101111111", "1000111101111110", "1000100101111111", "1001000101111101", "1001010001111011", "1000111001111101", "1000011101111111", "1000100101111111", "1000011101111111", "1001000101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100001111111", "1001100101111111", "1001100001111111", "1001100001111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001100001111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001111010000010", "1010000010000110", "1010000110000111", "1010001110000111", "1010001010000111", "1010000110000111", "1001111110000111", "1001101010000111", "1001011110000110", "1001011110000110", "1001010110000101", "1001010001111101", "1001001101111110", "1001001001111111", "1001001001111110", "1001001101111110", "1001001001111110", "1001001001111111", "1001011001111110", "1001111001111110", "1010000101111110", "1010000101111111", "1001111101111111", "1001111101111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000101111101", "1001101101111101", "1001100101111101", "1001100101111100", "1001110001111101", "1001101101111101", "1001010001111011", "1000110001111100", "1000100001111110", "1000110001111101", "1000110001111101", "1000010001111100", "1000001001111101", "0111111101111101", "0111111101111100", "0111110101111010", "0111111001111011", "1000000001111101", "1000001001111110", "1000000101111111", "0111111101111111", "0111111101111111", "1000000001111111", "1000011001111111", "1000100001111111", "1000110001111111", "1001000101111110", "1001010101111101", "1001010101111111", "1001011101111111", "1000011101111110", "1000010101111111", "1001000001111111", "1001100101111111", "1001001101111111", "1000110101111111", "1000011101111111", "1000011001111111", "1000110101111101", "1001001001111110", "1001100001111101", "1001110001111100", "1001111101111011", "1001111101111010", "1010000101111001", "1010000001111010", "1010000001111000", "1001111101111000", "1001110101111000", "1001110001111001", "1001101001111001", "1001101001111001", "1001101101111001", "1001110001111001", "1001110101111001", "1001111101111010", "1010000001111001", "1010000101111010", "1010000001111001", "1010000101111001", "1010000101111001", "1001111101110111", "1001000001111000", "1000010101111011", "1001010101111010", "1001100101111010", "1001110001111010", "1001110001111010", "1001101001111011", "1001011101111010", "1001010101111101", "1000100101111110", "1000100001111111", "1000110001111111", "1000111101111110", "1000100101111111", "1001000101111101", "1001010001111011", "1001000101111101", "1000011101111110", "1000100101111111", "1000100001111111", "1001010101111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001101001111111", "1001101001111111", "1001100101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100001111111", "1001011101111111", "1001100001111111", "1001100001111111", "1001011101111111", "1001100101111111", "1001100101111111", "1001110010000000", "1001111110000101", "1010000110000111", "1010001110000111", "1010001110000111", "1010000110000111", "1001111110000111", "1001100110000111", "1001011010000111", "1001010010000111", "1001011010000110", "1001011010000101", "1001010001111110", "1001001101111110", "1001001001111110", "1001001001111110", "1001000101111110", "1001000101111110", "1001001001111111", "1001011001111101", "1001111101111101", "1010000101111110", "1010000001111111", "1001111101111111", "1001111101111111", "1001111101111111", "1010000101111111", "1010001001111110", "1010000101111101", "1001101001111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001011001111100", "1001011001111100", "1000111101111110", "1000111001111110", "1000101101111100", "1000011001111101", "1000000101111101", "1000000001111101", "0111111001111011", "0111111001111011", "0111110001111010", "0111111001111010", "0111111101111100", "1000001001111110", "1000001001111110", "0111111101111111", "0111111101111111", "1000010101111110", "1001000101111110", "1001010101111101", "1001000001111110", "1001001101111100", "1001100001111101", "1001000101111111", "1001001101111111", "1000011101111111", "1000011001111110", "1001011101111111", "1001100101111111", "1001000101111111", "1000100001111111", "1000010001111111", "1000011001111110", "1000111001111101", "1001001001111101", "1001011101111101", "1001110001111011", "1001111101111010", "1010000001111010", "1010000101111001", "1010000001111010", "1010000101111001", "1010000001111000", "1001111001111000", "1001111101110111", "1001110001111000", "1001110001111000", "1001110001111001", "1001110101111000", "1001111101111000", "1010000001111001", "1010000001111010", "1001111101111010", "1001111101111010", "1001111101111010", "1010001001111001", "1001111101111000", "1001010001111000", "1000001101111011", "1001001101111010", "1001101001111010", "1001110001111010", "1001110001111010", "1001100101111011", "1001100001111011", "1001001001111101", "1000010001111110", "1000100001111111", "1000111001111111", "1000111101111110", "1000100101111111", "1001000101111101", "1001010001111011", "1001001001111101", "1000100001111111", "1000011101111111", "1000110001111111", "1001100001111111", "1001101001111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001101101111111", "1001111110000011", "1010000010000111", "1010001010000111", "1010001010000111", "1010000110001000", "1001111110001000", "1001100110000111", "1001010110000111", "1001010110000111", "1001010110000111", "1001010110000101", "1001010010000101", "1001010101111101", "1001010001111110", "1001001101111111", "1001001001111110", "1001000101111111", "1001000101111110", "1001000101111111", "1001010101111110", "1001111001111110", "1010000101111110", "1010000001111111", "1001111101111111", "1001111101111111", "1010000001111111", "1010000101111111", "1010001001111110", "1010000001111110", "1001101001111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001010101111101", "1001011101111011", "1000110101111101", "1000100101111101", "1000011101111101", "1000001001111100", "1000000101111101", "0111111101111100", "0111111101111011", "0111111001111100", "0111110101111011", "0111111101111010", "0111111101111101", "0111111101111111", "0111111101111111", "1000000101111111", "1000000101111111", "1000010001111110", "1000100101111110", "1001000101111110", "1001100101111101", "1001100001111110", "1001000101111110", "1000101101111111", "1000011001111111", "1000001101111110", "1000111101111111", "1001100101111111", "1001010101111111", "1000111101111111", "1000001101111111", "1000010101111111", "1000011101111110", "1000111101111101", "1001001001111101", "1001011101111101", "1001110001111011", "1001111001111011", "1001111101111010", "1010000101111001", "1010000101111001", "1010000101111010", "1010000001111001", "1010000001111000", "1010000001111000", "1001111101111000", "1001111001111000", "1001111101111000", "1001111101111000", "1001111101111001", "1001111101111010", "1001111101111010", "1001111101111010", "1010000101111001", "1010000001111010", "1010000101111010", "1010000001111000", "1001100101110111", "1000010001111011", "1001000101111010", "1001101101111010", "1001110001111010", "1001110001111010", "1001100101111010", "1001100001111011", "1000101001111110", "1000001101111110", "1000100001111111", "1000111101111111", "1000111101111110", "1000100101111111", "1001000001111101", "1001010001111011", "1001010001111100", "1000101101111111", "1000011101111111", "1001000101111111", "1001100101111111", "1001101101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001110010000001", "1001111110000111", "1010000110001000", "1010001010001000", "1010000110001000", "1001111110001001", "1001100110001000", "1001011010000111", "1001011010000111", "1001010110000111", "1001010010000110", "1001010010000101", "1001001110000101", "1001011001111101", "1001010101111101", "1001010001111110", "1001001101111110", "1001001001111111", "1001000101111111", "1001000101111111", "1001010001111110", "1001111001111110", "1010000101111110", "1010000101111111", "1001111101111111", "1001111101111111", "1001111101111111", "1010000101111111", "1010001001111110", "1010000101111110", "1001101001111101", "1001100101111101", "1001101001111101", "1001101101111100", "1001100101111101", "1001100101111101", "1000110001111110", "1000100101111101", "1000010001111100", "1000010001111101", "1000000001111101", "1000000001111101", "0111111101111100", "0111111101111100", "0111111101111100", "0111111101111001", "1000000001111101", "1000000001111110", "1000000101111111", "1000001101111110", "1000001001111111", "1000011101111111", "1000110001111111", "1001001001111111", "1001011001111111", "1001010001111111", "1000100001111111", "1000010001111110", "1000010001111110", "1000101001111111", "1001011101111110", "1001010101111101", "1001001101111101", "1001000101111110", "1000011001111110", "1000011001111111", "1000011001111110", "1000111101111101", "1001001001111101", "1001011101111100", "1001101101111100", "1001111001111011", "1001111101111010", "1010000101111010", "1010001001111000", "1010000101111010", "1010000101111001", "1010000001111000", "1010000001111001", "1010000001111000", "1001111101111000", "1001111101111000", "1001111101111001", "1001111101111010", "1001111101111010", "1001111101111010", "1010001001111001", "1010000101111001", "1010000101111010", "1010001101111001", "1010000101111001", "1001110001110111", "1000110001111011", "1001001001111011", "1001110001111010", "1001110101111010", "1001101001111011", "1001100101111010", "1001010001111101", "1000010001111111", "1000010001111101", "1000100101111110", "1000111001111111", "1000111101111110", "1000101001111111", "1000111001111110", "1001010001111010", "1001010101111011", "1000110101111110", "1000011101111111", "1001010001111111", "1001101101111111", "1001101001111111", "1001100101111111", "1001100001111111", "1001100001111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001101001111111", "1001111010000100", "1010000010001000", "1010000110001001", "1010000110001001", "1010000010001001", "1001101010001000", "1001011110000111", "1001011010000111", "1001011110000111", "1001011010000111", "1001010010000110", "1001001010000110", "1001001010000110", "1001011001111101", "1001011001111101", "1001010101111101", "1001010001111101", "1001001101111110", "1001001101111110", "1001001101111110", "1001010101111110", "1001111101111101", "1010000101111110", "1010000101111111", "1001111101111111", "1001111101111111", "1001111101111111", "1010000101111111", "1010001001111101", "1010000101111110", "1001101001111101", "1001100101111101", "1001101001111101", "1001110001111101", "1001101101111101", "1001010001111101", "1000110001111110", "1000100001111101", "1000011101111011", "1000010001111101", "1000000101111110", "0111111101111011", "1000000101111101", "0111111101111101", "0111111101111011", "0111111101111010", "1000000001111101", "1000000001111100", "1000001101111110", "1000010101111110", "1000011001111111", "0111111101111111", "1000010101111111", "1000011001111110", "1000110001111110", "1000110001111110", "1000010101111101", "1000011001111110", "1000001101111111", "1001000101111101", "1001001101111110", "1001001001111110", "1001000001111101", "1000100101111111", "1000010001111101", "1000011101111110", "1000011101111101", "1000111001111110", "1001001001111101", "1001011101111100", "1001101101111100", "1001110101111011", "1010000001111010", "1010000101111010", "1010001001111001", "1010000101111010", "1010000101111001", "1010000101111000", "1010000001111001", "1010000001111001", "1001111101111001", "1001111101111000", "1001111101111001", "1001111101111010", "1001111101111010", "1001111101111010", "1010000101111010", "1001100101111101", "1001111001111010", "1010000001111010", "1010001001111010", "1001111101111000", "1001010001111001", "1001011101111010", "1001110001111011", "1001110001111010", "1001101001111010", "1001100101111011", "1000101001111110", "1000000101111111", "1000010001111111", "1000101001111111", "1000111101111111", "1000111001111111", "1000101101111111", "1000110001111111", "1001010001111100", "1001010001111100", "1000111101111101", "1000101001111111", "1001011101111111", "1001110001111111", "1001100101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001110001111111", "1010000110000110", "1010000010001001", "1010000110001001", "1010000010001001", "1001101110001000", "1001100010001000", "1001011010000111", "1001010110000111", "1001010010000111", "1001010010000111", "1001001110000110", "1001001010000110", "1001001110000110", "1001011001111101", "1001010101111101", "1001010101111101", "1001010101111101", "1001010101111101", "1001001101111110", "1001010001111101", "1001011101111101", "1001111001111110", "1010000001111110", "1010000001111111", "1001111101111111", "1010000001111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000001111110", "1001101001111101", "1001100101111101", "1001101001111101", "1001110001111101", "1001110001111101", "1001010001111101", "1001000001111110", "1000011101111110", "1000100101111101", "1000001101111110", "1000000101111101", "1000000001111011", "0111111101111100", "0111111101111100", "0111111101111011", "0111111101111010", "1000000101111011", "1000000101111011", "1000000101111111", "1000100001111111", "1000110101111111", "1000010001111111", "0111111101111111", "1000010001111110", "1000101001111101", "1000100001111110", "1000100101111111", "1000100101111110", "1000110001111110", "1001010101111101", "1001010101111110", "1001000001111101", "1000011101111111", "1000010101111101", "1000010001111101", "1000011101111101", "1000011101111101", "1000111101111101", "1001001001111101", "1001011101111101", "1001110001111011", "1001111001111011", "1001111101111010", "1010000001111010", "1010001001111001", "1010000101111001", "1010000101111001", "1010000001111001", "1010000001111001", "1010000001111001", "1001111101111001", "1001111101111001", "1001111101111001", "1001111101111010", "1001111101111010", "1010000001111010", "1010000101111010", "1010000101111010", "1010001001111010", "1001111101111010", "1001111001111010", "1001101001111001", "1001010101111010", "1001100101111010", "1001101001111010", "1001101001111011", "1001100101111010", "1001010001111101", "1000010001111110", "1000000101111111", "1000010001111110", "1000101101111111", "1000111101111111", "1000111101111111", "1000110001111111", "1000100101111111", "1001001101111101", "1001010101111100", "1001000001111101", "1000111101111111", "1001101101111111", "1001110001111111", "1001100101111111", "1001100001111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100001111111", "1001011101111111", "1001100101111111", "1001111010000001", "1010000110000111", "1010000110001001", "1010000110001001", "1001110110001001", "1001100010001000", "1001011110000111", "1001011010000111", "1001010110000111", "1001001110000111", "1001001110000111", "1001001110000111", "1001001110000110", "1001001110000110", "1001010101111101", "1001010101111101", "1001010101111101", "1001010101111101", "1001010101111101", "1001010001111110", "1001011101111101", "1001100101111101", "1001111001111101", "1010000001111101", "1010000001111111", "1010000001111111", "1010000001111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000101111110", "1001101001111101", "1001100101111101", "1001100101111101", "1001110001111101", "1001110001111101", "1001011101111101", "1000100001111111", "1000010101111101", "1000010001111110", "1000001001111101", "1000001101111101", "1000000001111101", "0111111101111101", "0111111101111011", "0111111101111011", "0111111001111010", "1000000101111011", "1000000101111010", "1000010001111101", "1000100101111111", "1001010001111111", "1001010001111111", "1000000101111111", "1000011101111110", "1000110001111111", "1000111001111101", "1001010001111101", "1001001101111101", "1001010001111110", "1001100001111111", "1001000001111111", "1000011101111111", "1000011001111101", "1000011101111101", "1000011101111101", "1000100001111110", "1000100001111110", "1000111101111101", "1001001101111101", "1001011101111100", "1001110001111011", "1001111001111011", "1001111101111010", "1010000101111010", "1010000101111001", "1010000101111001", "1010000001111010", "1010000001111010", "1010000101111001", "1010000001111010", "1010000001111001", "1001111101111000", "1001111101111000", "1001111101111001", "1010000001111001", "1010000001111001", "1010000001111010", "1010000101111001", "1001111101111001", "1001110101111010", "1001010001111010", "1000111101111010", "1001010101111010", "1001100101111010", "1001101001111010", "1001101001111011", "1001100001111100", "1000100101111101", "1000001001111111", "1000000001111111", "1000010101111110", "1000110001111111", "1000111101111111", "1000111101111111", "1000110101111111", "1000101101111111", "1001000101111101", "1001010101111011", "1001001101111100", "1001001101111110", "1001110001111111", "1001110001111111", "1001100101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100101111111", "1001111110000011", "1010000110000111", "1010000110001001", "1001111110001001", "1001100110000111", "1001011110001000", "1001011010000111", "1001010110000111", "1001010110000111", "1001010010000111", "1001010010000111", "1001010010000111", "1001001110000110", "1001000110000101", "1001010001111101", "1001010001111101", "1001010001111101", "1001010101111101", "1001010101111101", "1001010101111101", "1001011101111101", "1001100101111101", "1001110101111101", "1001111101111101", "1010000001111111", "1010000001111111", "1010000001111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000101111110", "1001101101111101", "1001100101111100", "1001101001111101", "1001110001111101", "1001111001111100", "1001011001111101", "1000100101111110", "1000011001111101", "1000010001111101", "1000001001111100", "1000000101111110", "1000000101111110", "1000000101111101", "0111111101111100", "0111111101111100", "0111111101111010", "1000000001111100", "1000000101111010", "1000010101111100", "1000101001111110", "1000111101111110", "1000111101111111", "1000100101111110", "1000011001111110", "1000111101111111", "1001010101111101", "1001001101111101", "1001000001111101", "1001011101111111", "1001010001111111", "1000100001111111", "1000011101111111", "1000011001111110", "1000011101111101", "1000011101111111", "1000100001111111", "1000100101111111", "1000111001111110", "1001001101111101", "1001011101111101", "1001101001111011", "1001111001111011", "1001111101111010", "1001111101111010", "1010000101111010", "1010000101111001", "1010000101111010", "1010000001111010", "1010000101111010", "1010000001111001", "1010000001111000", "1010000001111000", "1001111101111001", "1001111101111001", "1001111101111001", "1001111101111001", "1001111101111010", "1001111001111010", "1001010101111011", "1001011001111010", "1001010001111011", "1000111101111011", "1001010101111010", "1001100101111010", "1001101001111010", "1001100101111100", "1001001001111101", "1000001001111110", "1000000101111111", "1000000101111111", "1000100001111110", "1000110101111111", "1000111101111111", "1000111101111110", "1000111001111111", "1000101101111111", "1001000001111101", "1001010101111011", "1001010001111100", "1001100001111110", "1001110101111111", "1001101101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100001111111", "1001101001111111", "1010000010000100", "1010000110001000", "1010000010001001", "1001110010001001", "1001100010001001", "1001011110001000", "1001011110001000", "1001011110000111", "1001011010000111", "1001010110000111", "1001001110000111", "1001001010000110", "1001001010000110", "1001000110000101", "1001010001111110", "1001010001111110", "1001010001111110", "1001010001111101", "1001010001111101", "1001010101111101", "1001011001111101", "1001100101111101", "1001110001111101", "1001111001111110", "1010000001111111", "1010000001111111", "1010000101111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000101111101", "1001101101111101", "1001100101111100", "1001101001111101", "1001110001111101", "1001100101111101", "1001001101111101", "1000100101111111", "1000011101111101", "1000010001111101", "1000001001111110", "1000000101111110", "1000000101111110", "1000001101111110", "1000000101111101", "1000000101111101", "0111111101111100", "1000000001111100", "1000000101111010", "1000010101111010", "1000101101111110", "1000111001111101", "1000100101111111", "1000101101111110", "1001000101111110", "1001001101111101", "1001001101111101", "1000110101111110", "1001010101111111", "1001011101111111", "1000110101111111", "1000011001111111", "1000100001111111", "1000011101111101", "1000011101111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000111001111101", "1001001001111101", "1001010101111101", "1001101001111011", "1001110101111011", "1001111101111010", "1001111101111010", "1010000001111010", "1010000001111010", "1010000101111010", "1010000101111010", "1010000001111010", "1010000001111010", "1010000001111001", "1010000001111001", "1001111101111001", "1001111101111010", "1001111101111010", "1001111001111010", "1001110001111010", "1001110001111001", "1000111101111010", "1001000001111010", "1001001101111010", "1000111101111011", "1001010101111010", "1001100101111011", "1001100101111011", "1001100001111101", "1000011101111111", "1000000101111111", "1000001001111110", "1000000101111111", "1000101001111110", "1000111001111111", "1000111101111110", "1000111101111111", "1000111001111111", "1000101101111111", "1000111101111110", "1001010101111011", "1001010001111101", "1001101101111110", "1001110101111111", "1001101101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100001111111", "1001101101111111", "1010000010000100", "1010000110001001", "1001111010001001", "1001100110001001", "1001011110001001", "1001011110001001", "1001011110001000", "1001011010000111", "1001011010000111", "1001010010000111", "1001000110000110", "1001001110000111", "1001001010000110", "1001000110000101", "1001001101111110", "1001001101111110", "1001001101111110", "1001001101111111", "1001010001111110", "1001010001111110", "1001011101111101", "1001100101111101", "1001101101111101", "1001111001111110", "1001111101111111", "1010000001111111", "1010000001111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000101111101", "1001101101111101", "1001100101111101", "1001101001111101", "1001100101111101", "1001101101111101", "1001000001111101", "1000101001111101", "1000010001111100", "1000001101111101", "1000001101111111", "1000001001111110", "1000000101111101", "1000001101111101", "1000010001111101", "1000000101111101", "1000000101111101", "1000000101111101", "1000001101111011", "1000001001111010", "1000111001111100", "1000100101111111", "1000110001111111", "1001011101111101", "1001010101111101", "1001010001111101", "1000111101111101", "1001001101111111", "1001011101111111", "1001000001111111", "1000010101111111", "1000011101111110", "1000110001111111", "1000011101111110", "1000100001111111", "1000100101111111", "1000101101111111", "1000100101111111", "1000110101111110", "1001001001111101", "1001010001111101", "1001100101111100", "1001110101111011", "1001111101111011", "1001111101111010", "1001111101111010", "1010000001111010", "1010000101111010", "1010000001111010", "1010000001111010", "1010000101111010", "1010000001111010", "1001111101111010", "1001111101111010", "1001111001111010", "1001111001111011", "1001111001111010", "1001110001111001", "1001110001111000", "1001010101111000", "1001000101111001", "1001001001111000", "1001010001110111", "1001011001111001", "1001100001111100", "1001100101111101", "1001001001111101", "0111111101111111", "1000001001111110", "1000001001111110", "1000010001111110", "1000101101111111", "1000111101111111", "1000111101111110", "1000111101111110", "1000111101111111", "1000110001111111", "1000111001111111", "1001010101111011", "1001011001111101", "1001110001111110", "1001110101111111", "1001100101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001110001111111", "1010000110000101", "1001111110001001", "1001100110001001", "1001011110001001", "1001011110001001", "1001011110001001", "1001011010000111", "1001011110001000", "1001011010000111", "1001001110000111", "1001000110000110", "1001000110000110", "1001000110000110", "1001000110000101", "1001000001111111", "1001000101111110", "1001001001111101", "1001001001111111", "1001001101111110", "1001010001111101", "1001011101111101", "1001100001111101", "1001110001111101", "1001111001111101", "1001111101111111", "1001111101111111", "1001111101111111", "1001111110000000", "1010000001111111", "1010001001111110", "1010000101111101", "1001101101111101", "1001100101111100", "1001100101111101", "1001101001111101", "1001110001111100", "1000111101111101", "1000011001111110", "1000010001111101", "1000010001111101", "1000010001111101", "1000000101111110", "1000000001111100", "1000000101111011", "1000001101111101", "1000000101111101", "1000000001111101", "1000001001111100", "1000001001111101", "1000001001111011", "1000010001111010", "1000011101111101", "1001100001111101", "1000111101111100", "1000110001111110", "1000110001111111", "1001001101111110", "1001100101111111", "1001010001111110", "1000011101111111", "1000011101111101", "1000011101111110", "1000110001111110", "1000011101111110", "1000100101111111", "1000100101111111", "1000101101111111", "1000100101111111", "1000110001111111", "1001000001111101", "1001001101111101", "1001100101111100", "1001110001111011", "1001111001111011", "1001111001111011", "1001111101111010", "1001111101111010", "1010000001111010", "1010000001111010", "1010000001111010", "1001111101111010", "1001110001111011", "1001110101111011", "1001110101111011", "1001111001111010", "1001111101111010", "1001111101111010", "1001111101111001", "1001111101111010", "1001111101111001", "1001111101110111", "1001110001110111", "1001101001111001", "1001100101111010", "1001100101111101", "1001100001111100", "1000011001111111", "0111111101111111", "1000001001111110", "1000010001111101", "1000011101111110", "1000110001111111", "1000111001111111", "1000111101111110", "1000111101111110", "1000111101111110", "1000110001111111", "1000111001111111", "1001010101111011", "1001011101111101", "1001110101111110", "1001110101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001011101111111", "1001100001111111", "1001110001111111", "1010000010000110", "1001101110001000", "1001011110001001", "1001011010001001", "1001011110001001", "1001011110001001", "1001011010001000", "1001011010000111", "1001010010000111", "1001001010000111", "1001000110000111", "1001000010000110", "1001000110000110", "1001000110000101", "1000111001111111", "1000111101111111", "1001000001111111", "1001000101111111", "1001001101111110", "1001010001111101", "1001011101111101", "1001100101111101", "1001110001111101", "1001111101111110", "1010000001111111", "1001111101111111", "1001111101111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000101111101", "1001101101111101", "1001100101111101", "1001100101111101", "1001110001111101", "1001101001111100", "1000110101111110", "1000011101111110", "1000010001111110", "1000010001111110", "1000001001111110", "1000001001111101", "1000000101111101", "0111111101111010", "0111111101111010", "0111111101111100", "1000001001111100", "1000001001111101", "1000010001111011", "1000001101111101", "1000001001111101", "1000111001111101", "1001100101111011", "1001100101111101", "1000100101111111", "1000110001111101", "1001100101111110", "1001011101111111", "1000101001111111", "1000011101111110", "1000100101111111", "1000010001111110", "1000101001111111", "1000011001111101", "1000100001111111", "1000100101111111", "1000101101111111", "1000100101111110", "1000101101111111", "1000111101111110", "1001000101111101", "1001011101111100", "1001110001111011", "1001110101111011", "1001111101111010", "1001111101111010", "1001111101111010", "1001111101111010", "1001111101111010", "1001111101111010", "1001111101111010", "1001110001111011", "1001100101111100", "1001011101111100", "1001100101111011", "1001110001111010", "1001110001111010", "1001110001111010", "1001110101111001", "1001111101111000", "1001110101110111", "1001101101110111", "1001100001111010", "1001100101111101", "1001101001111101", "1001001001111101", "0111111101111111", "1000000001111111", "1000010001111101", "1000010001111101", "1000100101111110", "1000110001111111", "1000111101111111", "1001000001111110", "1000111101111111", "1000111101111111", "1000110001111111", "1000110101111111", "1001010101111011", "1001100101111101", "1001110101111110", "1001110001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001111010000001", "1001111110000111", "1001100110001001", "1001010110001000", "1001011010001000", "1001011010001000", "1001011010001000", "1001010110001000", "1001010110000111", "1001010010000111", "1001001010000111", "1001000110000111", "1001000110000110", "1001001010000111", "1001001010000110", "1000110101111111", "1000110101111111", "1000111101111111", "1001000101111111", "1001010001111101", "1001010001111101", "1001011101111101", "1001101001111101", "1001110101111101", "1001111101111101", "1001111101111111", "1001111101111111", "1001111110000000", "1001111110000000", "1010000101111111", "1010001001111101", "1010000001111110", "1001101001111101", "1001100101111100", "1001100101111101", "1001101101111101", "1001100001111101", "1000111001111101", "1000011101111111", "1000010001111101", "1000001001111110", "1000000101111110", "1000001101111110", "1000001001111101", "0111111101111010", "0111111101111011", "0111111101111100", "0111111101111011", "1000010001111100", "1000010101111101", "1000100001111101", "1000010101111100", "1001000101111010", "1010011101111110", "1010000101111101", "1000100101111110", "1001011101111110", "1001101101111111", "1001000101111110", "1000001001111111", "1000100001111110", "1000011101111101", "1000000101111111", "1000100001111111", "1000011101111101", "1000100001111111", "1000100101111111", "1000101001111111", "1000100101111110", "1000101101111111", "1000111001111110", "1001000001111101", "1001011001111101", "1001101101111011", "1001110101111011", "1001111001111010", "1001111001111011", "1001111001111010", "1001111001111010", "1001111001111010", "1001111101111010", "1010000001111010", "1010000101111010", "1010000001111010", "1001111101111010", "1010000001111001", "1010000101111000", "1010001001110110", "1001111001110100", "1001100101110011", "1001100101110010", "1001010001110100", "1001100101110101", "1001100101111001", "1001100101111100", "1001011101111101", "1000010001111111", "0111111101111111", "1000001101111110", "1000010001111110", "1000010101111110", "1000100101111111", "1000101001111111", "1000111101111111", "1001000001111110", "1000111101111110", "1000111101111111", "1000111001111111", "1000111001111111", "1001010001111011", "1001100101111101", "1001111001111110", "1001101101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001110110000001", "1001110010000111", "1001011010001000", "1001011010001000", "1001011010001000", "1001010110001001", "1001010010001000", "1001010010001000", "1001010010001000", "1001001110000111", "1001001110000111", "1001001110000111", "1001001110000111", "1001010010000111", "1001010010000111", "1000110001111111", "1000111001111110", "1000111101111111", "1001000101111110", "1001001101111111", "1001010001111110", "1001011101111101", "1001101001111101", "1001110101111101", "1010000001111101", "1010000101111111", "1001111101111111", "1001111110000000", "1001111110000000", "1010000101111111", "1001111101111101", "1001110001111101", "1001101001111101", "1001100001111101", "1001101001111101", "1001100101111101", "1001011101111101", "1000101101111110", "1000010101111100", "1000010101111101", "1000010001111101", "1000000101111101", "1000010001111101", "1000001101111101", "0111111101111010", "0111111101111010", "1000000101111101", "1000000001111100", "1000000101111011", "1000010001111100", "1000010001111101", "1000011001111010", "1001001101111010", "1010000101111101", "1001011101111110", "1001000101111110", "1001110101111111", "1001100101111111", "1000011101111111", "1000001001111110", "1000011001111101", "1000011101111100", "1000000101111111", "1000010101111101", "1000011101111101", "1000011101111101", "1000100101111111", "1000101001111111", "1000101001111111", "1000100101111111", "1000111001111110", "1000111001111110", "1001010001111101", "1001100101111100", "1001110001111100", "1001111001111011", "1001111001111010", "1001111001111011", "1001110101111011", "1001111001111011", "1001111101111010", "1010000001111010", "1010000101111010", "1010000001111010", "1001111101111011", "1001111101111010", "1010000001111010", "1010001001111000", "1010000101110110", "1001111101110101", "1001111101110101", "1001111101110101", "1001101001111000", "1001100001111011", "1001011101111100", "1000111101111110", "0111111101111111", "0111111101111111", "1000010001111111", "1000011001111101", "1000011101111110", "1000101001111111", "1000101101111111", "1001000001111110", "1001000101111101", "1000111101111110", "1000111101111110", "1000111101111110", "1000111101111110", "1001010001111100", "1001100101111100", "1001111001111110", "1001100101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001110110000001", "1001100110001000", "1001010010001000", "1001010110001000", "1001010110000111", "1001010010001000", "1001010010001000", "1001001110001000", "1001001110001000", "1001001110000111", "1001010010000111", "1001011010000111", "1001011110000111", "1001011110000111", "1001011110000111", "1000101001111111", "1000101101111111", "1000111001111111", "1001000001111110", "1001000101111111", "1001001101111110", "1001011101111101", "1001100101111110", "1001111001111101", "1010000101111101", "1010000101111111", "1001111101111111", "1001111101111111", "1001111110000000", "1010000101111111", "1010001101111101", "1010000101111101", "1001101001111101", "1001100001111101", "1001101001111101", "1001100101111101", "1001010001111101", "1000100101111111", "1000011101111011", "1000011001111101", "1000010001111110", "1000000101111101", "1000010001111101", "1000001001111101", "0111111101111001", "0111111101111011", "0111111101111010", "1000000001111010", "1000001001111110", "1000000001111010", "1000001001111001", "1000111001111100", "1001000101111100", "1001011101111011", "1000111101111101", "1001100101111111", "1001100110000001", "1000110001111111", "1000001001111110", "1000000101111111", "1000011001111101", "1000011101111100", "1000000101111111", "1000011001111101", "1000010001111101", "1000011101111101", "1000100101111110", "1000100101111111", "1000101001111111", "1000100101111111", "1000110001111111", "1000110101111111", "1001000101111110", "1001011101111100", "1001101101111100", "1001110101111011", "1001110101111100", "1001110001111100", "1001111001111100", "1001111001111010", "1001111001111011", "1001111101111010", "1001111101111010", "1001111101111010", "1001111101111011", "1001111001111011", "1001111001111011", "1001111001111011", "1001111101111010", "1001111001111010", "1001110101111010", "1001101101111011", "1001011101111100", "1001100101111100", "1001001001111101", "1000100101111110", "0111111101111111", "0111111101111111", "1000011001111101", "1000011101111110", "1000100101111111", "1000101101111111", "1000110001111111", "1001000101111110", "1001000101111101", "1000111101111110", "1001000001111110", "1001000001111110", "1000111101111111", "1001010001111011", "1001100101111101", "1001110001111101", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001110010000010", "1001011010000111", "1001001110001001", "1001010010001000", "1001010010001000", "1001010010001000", "1001001010000111", "1001001010001000", "1001010110001000", "1001011010001000", "1001011110001000", "1001011110000111", "1001011110000111", "1001011010000111", "1001011010001000", "1000100101111111", "1000101001111111", "1000110001111111", "1000111101111111", "1001000001111111", "1001010001111101", "1001100101111101", "1001101001111101", "1001111001111101", "1010000101111101", "1010000101111111", "1001111101111111", "1010000001111111", "1010000001111111", "1010000101111111", "1010001101111101", "1010000101111101", "1001101001111101", "1001011101111101", "1001100001111101", "1001100001111101", "1000110001111110", "1000011101111111", "1000100001111101", "1000011001111110", "1000000001111111", "1000001101111101", "1000010001111110", "1000001001111101", "0111111101111000", "1000000001111010", "0111111101111010", "1000000001111010", "1000000101111010", "1000000101111011", "1000001001111001", "1000111101111100", "1000101101111010", "1001000101111011", "1000111001111101", "1001110010000001", "1001000101111111", "1000001001111111", "1000000101111111", "0111111101111111", "1000011101111101", "1000011101111101", "1000000101111111", "1000011001111101", "1000010001111101", "1000010101111101", "1000100001111110", "1000100101111111", "1000101001111111", "1000100001111111", "1000101101111111", "1000110001111111", "1000110001111111", "1001010001111101", "1001100001111101", "1001101101111100", "1001110001111100", "1001110001111100", "1001110101111011", "1001110101111100", "1001111001111011", "1001111001111011", "1001111101111010", "1001111101111010", "1001111101111010", "1001111101111010", "1001111001111011", "1001111001111010", "1001110101111010", "1001111001111010", "1001110001111010", "1001100101111100", "1001100001111100", "1001011101111100", "1000101101111101", "1000011101111110", "0111111101111111", "1000000101111111", "1000011101111110", "1000011101111111", "1000011101111111", "1000101001111111", "1000101001111111", "1001001001111101", "1001000101111110", "1001000001111110", "1001000001111110", "1001000101111101", "1000111101111110", "1001001101111100", "1001100101111100", "1001110001111101", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001010101111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001101110000010", "1001010010000111", "1001001110001001", "1001010010001000", "1001001010001001", "1001001110001000", "1001010010001000", "1001010010001000", "1001011010001000", "1001011010001000", "1001010110001000", "1001011110000111", "1001010110000111", "1001010110000111", "1001011010000111", "1000100101111111", "1000100101111111", "1000101001111111", "1000110101111111", "1000111101111111", "1001010101111101", "1001101001111101", "1001110001111101", "1001111001111110", "1010000101111101", "1010000101111110", "1001111101111111", "1001111110000000", "1001111110000000", "1010000001111111", "1010001101111110", "1010000101111101", "1001101101111101", "1001011101111101", "1001011101111101", "1001011001111101", "1000111001111110", "1000101101111110", "1000011101111110", "1000010001111110", "0111111101111111", "1000001101111111", "1000010001111111", "1000001101111101", "0111111101111010", "0111111101111010", "0111111101111010", "0111111101111010", "1000000001111010", "1000001001111100", "1000000101111010", "1001100001111010", "1001000101111010", "1001000101111101", "1000111101111110", "1001000101111111", "1000011101111110", "1000000101111111", "0111111101111111", "1000000001111111", "1000011101111101", "1000011101111101", "1000001001111110", "1000011001111101", "1000011001111101", "1000010001111101", "1000011001111110", "1000100001111111", "1000101001111111", "1000100001111110", "1000101001111111", "1000101001111111", "1000100101111111", "1000111001111111", "1001001001111101", "1001011101111101", "1001100101111100", "1001101101111100", "1001110001111100", "1001110101111011", "1001110101111010", "1001111001111010", "1001110101111011", "1001110101111011", "1001110101111010", "1001110001111010", "1001110101111010", "1001110001111001", "1001101001111001", "1001101001111001", "1001101101111001", "1001101001111010", "1001011101111100", "1001000101111101", "1000100001111110", "1000010001111111", "1000000101111111", "1000001001111110", "1000100001111110", "1000100101111111", "1000100101111111", "1000100101111111", "1000110101111111", "1001001001111101", "1001000101111101", "1001000001111110", "1001000101111101", "1001000101111110", "1001000001111110", "1001001101111100", "1001100101111100", "1001101001111101", "1001011101111111", "1001011001111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001010101111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001010101111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001100110000011", "1001001110001000", "1001000110001001", "1001001110001001", "1001010010001000", "1001010010001001", "1001010010001000", "1001010010001000", "1001010010001001", "1001010010001000", "1001010110000111", "1001011010000111", "1001011110000111", "1001100010000110", "1001100110000101", "1000100101111111", "1000100101111111", "1000100101111111", "1000101101111111", "1000110101111111", "1001011001111101", "1001101001111101", "1001101101111110", "1001111001111101", "1010000101111101", "1010000101111111", "1001111101111111", "1001111101111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000101111101", "1001101001111101", "1001011101111101", "1001011101111101", "1001010001111101", "1000101101111111", "1000100101111110", "1000010101111110", "1000010101111101", "1000000001111111", "1000001001111111", "1000010001111110", "1000010001111110", "1000000101111011", "0111111101111101", "0111111101111100", "0111111101111010", "0111111101111001", "1000000101111010", "1000001001111011", "1001000101111001", "1001100101111010", "1000111001111110", "1000111101111110", "1000100101111110", "1000010101111110", "1000001001111111", "1000001001111110", "1000001101111110", "1000100101111110", "1000011101111101", "1000010001111101", "1000011001111110", "1000010001111110", "1000010001111110", "1000010001111101", "1000011101111101", "1000100001111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000101101111111", "1000100001111110", "1000111001111111", "1001010001111101", "1001011101111101", "1001101001111100", "1001110001111100", "1001110001111100", "1001110101111010", "1001110101111010", "1001110001111010", "1001110001111010", "1001101001111001", "1001101101111000", "1001101101111000", "1001101001111001", "1001100101111001", "1001100101111001", "1001100101111010", "1001011101111011", "1000110101111110", "1000101101111110", "1000001101111111", "1000000101111111", "1000001101111110", "1000100101111110", "1000100101111111", "1000100101111111", "1000100101111111", "1000111101111111", "1001001101111101", "1001001001111101", "1001000101111101", "1001001001111101", "1001001001111101", "1001000001111110", "1001001101111100", "1001100101111100", "1001100001111110", "1001011001111111", "1001011001111111", "1001011101111111", "1001010101111111", "1001010101111111", "1001010001111111", "1001010001111111", "1001010101111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001011001111111", "1001010001111111", "1001011001111111", "1001011001111111", "1001011101111111", "1001100010000100", "1001000110001000", "1001001010001000", "1001011010001001", "1001011010001001", "1001011010001000", "1001010010001000", "1001010010001000", "1001010010000111", "1001011110000111", "1001011110000110", "1001100110000101", "1001100110000101", "1001100110000100", "1001101110000011", "1000100101111111", "1000100101111110", "1000100101111111", "1000100101111111", "1000110001111111", "1001010001111101", "1001100101111101", "1001101101111101", "1001111001111110", "1010000101111101", "1010000001111111", "1001111101111111", "1010000001111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000101111101", "1001101001111101", "1001011101111101", "1001100001111101", "1000110101111111", "1000100001111111", "1000011101111101", "1000011101111110", "1000011001111110", "1000001101111111", "1000001101111110", "1000001001111110", "1000001001111110", "1000000101111010", "1000001101111101", "1000001001111101", "1000000101111100", "1000000001111010", "1000000001111000", "0111111101111000", "1000100001111001", "1001000001111011", "1000111101111110", "1000110101111111", "1000100001111110", "1000000101111111", "1000000001111111", "1000000101111111", "1000001101111110", "1000100101111111", "1000100101111110", "1000010001111101", "1000011101111110", "1000010001111101", "1000011001111101", "1000010001111101", "1000010001111101", "1000100001111110", "1000100001111110", "1000011101111110", "1000100101111111", "1000100101111111", "1000101101111111", "1000100101111110", "1000010001111101", "1000101001111111", "1001000101111110", "1001011001111101", "1001100101111101", "1001101101111100", "1001110001111011", "1001110001111010", "1001111001111010", "1001110101111010", "1001110101111001", "1001110001111000", "1001101001111000", "1001101001110111", "1001101001111000", "1001100101111010", "1001100101111011", "1001011101111100", "1000111001111111", "1000101101111111", "1000010001111101", "1000000001111111", "1000010101111101", "1000100101111111", "1000100001111111", "1000100101111111", "1000101001111111", "1000111101111111", "1001001101111101", "1001000101111101", "1001000101111101", "1001001001111101", "1001001001111101", "1001000001111110", "1001010001111100", "1001101001111101", "1001011101111110", "1001011101111111", "1001011001111111", "1001010101111111", "1001010101111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001010101111111", "1001010101111111", "1001011001111111", "1001011101111111", "1001100010000101", "1001000110001000", "1001010010001001", "1001011110001001", "1001011110001001", "1001010110001000", "1001010110001000", "1001011010000111", "1001011110000110", "1001100010000101", "1001101010000101", "1001110010000100", "1001111010000001", "1001110001111111", "1001100001111111", "1000100101111111", "1000100001111101", "1000100001111111", "1000100101111111", "1000101001111111", "1001000101111110", "1001011101111101", "1001101001111110", "1001111001111110", "1010000101111101", "1010000101111111", "1001111101111111", "1001111101111111", "1010000001111111", "1010000101111111", "1010001101111101", "1010000001111101", "1001101001111101", "1001011101111111", "1001010101111110", "1001000001111110", "1000011101111101", "1000100101111111", "1000100101111111", "1000011101111111", "1000010101111110", "1000001101111110", "1000000101111111", "1000000101111111", "1000000001111010", "1000000101111010", "1000010001111101", "1000001001111101", "1000010001111010", "1000000101111010", "0111111101111010", "1000000001111001", "1000011101111001", "1000100001111010", "1000110001111100", "1000011001111110", "1000000101111111", "0111111101111111", "1000000101111111", "1000010001111101", "1000110001111111", "1000100101111110", "1000010001111110", "1000100001111110", "1000010001111101", "1000010101111101", "1000010001111101", "1000010001111101", "1000011001111101", "1000011101111111", "1000100101111111", "1000100101111111", "1000101001111111", "1000101001111111", "1000110101111111", "1000110001111111", "1000101001111111", "1000111001111111", "1001000101111111", "1001001101111110", "1001011001111101", "1001011101111101", "1001100101111100", "1001110001111011", "1001101101111010", "1001110001111010", "1001110001111000", "1001101001111000", "1001100101111001", "1001101101111001", "1001100101111010", "1001011101111011", "1001101001111101", "1000110101111111", "1000100001111111", "1000010001111111", "1000000101111111", "1000011101111110", "1000100101111111", "1000100101111111", "1000100101111111", "1000101001111111", "1000111101111110", "1001001101111101", "1001001001111101", "1001000101111110", "1001001101111101", "1001001001111101", "1001000101111101", "1001010001111100", "1001101101111101", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001010001111111", "1001010101111110", "1001010001111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001010101111111", "1001010101111110", "1001010101111111", "1001010101111111", "1001011110000000", "1001011110000111", "1001010010001001", "1001011110001001", "1001011110001001", "1001011110001000", "1001011110000111", "1001100010000111", "1001100110000101", "1001101110000100", "1001110010000010", "1001111010000001", "1001101101111111", "1001010001111111", "1000111101111111", "1000111101111111", "1000101101111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000111101111111", "1001010101111110", "1001100001111110", "1001110101111110", "1010000001111101", "1010000001111111", "1001111101111111", "1001111101111111", "1010000101111111", "1010000101111111", "1010001101111101", "1010000001111110", "1001011101111111", "1001000101111111", "1001001001111110", "1000111101111111", "1000010001111110", "1000100001111111", "1000011101111110", "1000011101111111", "1000011001111110", "1000010001111110", "1000001001111110", "1000010001111101", "1000001101111010", "1000000101111010", "1000010001111100", "1000010001111101", "1000010001111101", "1000000001111100", "0111111101111000", "0111111101111010", "1000000001111000", "1000011001111010", "1000101001111101", "1000100001111010", "1000011101111101", "1000000101111111", "1000001101111110", "1000011101111101", "1000111101111111", "1000100101111101", "1000010001111110", "1000100101111101", "1000010001111101", "1000010001111101", "1000010001111101", "1000010101111101", "1000010001111101", "1000011001111101", "1000100001111110", "1000100101111111", "1000100101111111", "1000100101111111", "1000111001111111", "1001000101111101", "1001010001111101", "1001011101111101", "1001100101111100", "1001101101111011", "1001100101111100", "1001100101111011", "1001100101111100", "1001100101111011", "1001100101111100", "1001101001111011", "1001101001111011", "1001101001111010", "1001100101111010", "1001100101111010", "1001011101111010", "1001010001111010", "1001001101111101", "1001000101111101", "1000110001111111", "1000010001111111", "1000010001111110", "1000011101111111", "1000100101111111", "1000100101111111", "1000100001111110", "1000101101111111", "1001000001111110", "1001001101111101", "1001001001111101", "1001000101111101", "1001010001111101", "1001010001111101", "1001000101111101", "1001011001111100", "1001101101111101", "1001011101111111", "1001100101111111", "1001100101111111", "1001100101111110", "1001100101111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001010101111111", "1001010101111111", "1001010101111111", "1001010101111111", "1001010101111111", "1001010101111111", "1001010001111111", "1001010101111111", "1001100010000001", "1001010110000111", "1001011110001000", "1001100110000111", "1001011110000111", "1001011110000110", "1001100110000110", "1001101110000110", "1001110010000101", "1001110010000001", "1001110001111111", "1001100001111111", "1001000001111111", "1000111001111111", "1001001001111111", "1001010101111110", "1000110101111111", "1000110001111111", "1000101101111111", "1000101101111111", "1000101001111111", "1000111101111111", "1001010001111110", "1001011101111101", "1001110001111110", "1010000101111101", "1010000101111110", "1001111101111111", "1010000001111111", "1010000001111111", "1010000101111111", "1010001001111101", "1001101001111111", "1001010101111111", "1001010101111110", "1000111101111111", "1000100101111110", "1000000001111111", "1000011101111111", "1000100101111111", "1000011101111111", "1000011001111101", "1000011101111101", "1000010001111110", "1000010101111101", "1000001001111100", "1000010001111010", "1000000101111010", "1000001101111101", "1000010001111101", "1000000101111010", "0111111101111010", "0111111101111010", "0111111101111010", "1000011001111010", "1000100001111101", "1000110001111111", "1000011101111010", "1000010001111011", "1000010101111101", "1000101001111111", "1000111101111111", "1000100101111110", "1000010101111110", "1000100101111110", "1000010101111101", "1000001001111110", "1000010101111101", "1000010001111101", "1000010101111101", "1000010101111101", "1000100001111110", "1000100101111111", "1000101001111111", "1000101001111111", "1000110101111111", "1001000101111110", "1001011101111101", "1001101001111101", "1001101101111101", "1001101101111101", "1001101101111100", "1001101101111100", "1001101001111100", "1001101001111100", "1001110001111100", "1001110001111100", "1001110001111100", "1001110001111100", "1001110001111011", "1001110001111010", "1001100101111011", "1001011001111101", "1001000101111101", "1000111101111101", "1001000001111101", "1000111101111101", "1000110001111111", "1000100101111111", "1000100101111111", "1000100101111111", "1000011101111111", "1000110001111111", "1001000101111110", "1001010001111101", "1001000101111110", "1001000101111101", "1001001101111101", "1001001101111101", "1001000101111101", "1001011101111100", "1001101101111101", "1001100001111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001101001111110", "1001100101111111", "1001100001111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001010101111111", "1001010101111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001100110000001", "1001011110000111", "1001101110000111", "1001110010000110", "1001100010000110", "1001011110000101", "1001100110000101", "1001110010000100", "1001110110000001", "1001110101111111", "1001100101111111", "1001001101111111", "1001001001111111", "1001010101111101", "1001100001111101", "1001011101111101", "1000110001111101", "1000110101111110", "1000111001111111", "1000111001111111", "1000110101111111", "1001000001111111", "1001001001111110", "1001010001111110", "1001101001111110", "1010000001111101", "1010000101111110", "1010000001111111", "1010000101111111", "1010000101111111", "1001111001111111", "1001110101111110", "1001111001111110", "1001100101111110", "1001010001111101", "1001001101111110", "1000010001111110", "0111111101111111", "1000010001111111", "1000100001111111", "1000010101111111", "1000010001111110", "1000011101111101", "1000011001111110", "1000010001111110", "1000000101111110", "1000010001111011", "1000010101111100", "1000000101111100", "1000001001111010", "0111111101111010", "0111111101111100", "1000000001111100", "0111111101111010", "1000000101111010", "1000010001111011", "1000100101111010", "1000110001111101", "1000010001111011", "1000011101111100", "1000110001111111", "1001000001111111", "1000011101111101", "1000010101111110", "1000101101111101", "1000011001111101", "1000001101111110", "1000010001111101", "1000010101111101", "1000010001111101", "1000010101111101", "1000011101111101", "1000100101111111", "1000101001111111", "1000101001111111", "1000110001111111", "1001001001111101", "1001011101111101", "1001100101111101", "1001101101111101", "1001101101111101", "1001101101111101", "1001101001111100", "1001101001111011", "1001110101111011", "1001110101111011", "1001111001111011", "1001110101111011", "1001111001111011", "1001111001111011", "1001110001111100", "1001100001111100", "1001010101111101", "1001000101111101", "1001000101111101", "1001000001111110", "1000111101111110", "1000111101111101", "1000111101111101", "1000110101111110", "1000101001111111", "1000011101111111", "1000110001111111", "1001001001111110", "1001001101111110", "1001000101111101", "1001000101111101", "1001001101111110", "1001010001111101", "1001000101111101", "1001100101111101", "1001101001111110", "1001011101111111", "1001100101111111", "1001100001111111", "1001100001111111", "1001100001111111", "1001100101111111", "1001100101111111", "1001100001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111110", "1001011101111111", "1001011001111111", "1001010101111111", "1001101110000001", "1001101010000110", "1001110110001000", "1001101010000110", "1001100010000101", "1001100110000101", "1001101010000100", "1001101110000001", "1001110001111111", "1001011101111111", "1001010001111110", "1001011001111101", "1001011001111101", "1001011101111101", "1001100101111101", "1001100001111101", "1000100101111101", "1000101001111101", "1000110001111101", "1000111101111101", "1000111101111111", "1001000101111110", "1001000101111110", "1001000101111110", "1001100101111110", "1010000001111101", "1010000101111110", "1010000101111111", "1010000101111111", "1010000101111111", "1010000001111111", "1010001101111101", "1010000101111110", "1001100101111110", "1001010001111111", "1000101001111111", "1000001001111110", "0111111101111111", "1000000101111111", "1000011101111111", "1000010101111101", "1000000101111111", "1000011101111101", "1000011101111101", "1000010101111100", "1000010001111101", "1000010001111101", "1000010101111100", "1000010001111011", "1000001101111011", "1000000101111011", "0111111101111100", "1000000001111010", "1000010001111011", "0111111101111010", "1000010001111001", "1000110101111011", "1000100101111011", "1000101001111110", "1000100101111100", "1000110101111111", "1001000001111111", "1000011101111110", "1000011101111101", "1000101001111110", "1000011101111101", "1000010001111101", "1000001101111110", "1000011001111101", "1000010101111101", "1000010101111101", "1000011101111110", "1000100101111111", "1000110001111111", "1000101101111111", "1000110001111111", "1001001001111101", "1001011101111101", "1001100101111101", "1001101101111101", "1001110001111100", "1001110001111100", "1001101001111100", "1001110101111100", "1001111001111011", "1001111101111011", "1001111001111011", "1001111101111011", "1001111001111011", "1001110101111100", "1001101101111011", "1001100001111101", "1001010101111101", "1001001101111110", "1001001001111110", "1001000101111101", "1001000101111110", "1001000001111110", "1000111101111110", "1000110101111110", "1000110001111111", "1000100101111111", "1000110001111111", "1001001001111101", "1001010001111101", "1001000101111110", "1001000101111101", "1001001101111110", "1001010001111101", "1001000101111101", "1001101101111101", "1001100101111110", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001100001111111", "1001011101111111", "1001011001111111", "1001100001111111", "1001110001111111", "1001110001111111", "1001100101111111", "1001110110000010", "1001101110000111", "1001110010000111", "1001100110000110", "1001100110000101", "1001101110000100", "1001110110000001", "1001110101111111", "1001100001111111", "1001011001111110", "1001100001111110", "1001100001111101", "1001100001111101", "1001100101111101", "1001100101111101", "1001100001111101", "1000100101111110", "1000101001111101", "1000100101111101", "1000110001111101", "1000111101111110", "1001001001111110", "1001001001111111", "1001000101111110", "1001100101111110", "1010000001111110", "1010000101111101", "1010000101111111", "1010000001111111", "1010000101111111", "1010000101111111", "1010001101111101", "1001111101111111", "1001011101111110", "1001010101111101", "1000011001111110", "1000001101111110", "1000000101111111", "1000000001111111", "1000100101111101", "1000100101111101", "1000011101111101", "1000100101111011", "1000010101111110", "1000010001111101", "1000010001111101", "1000100001111101", "1000011001111110", "1000001001111101", "1000000101111100", "1000000001111101", "1000000001111101", "1000000101111100", "1000010001111010", "1000010001111001", "1000000101111000", "1000100101111100", "1000101001111101", "1000011101111011", "1000101001111101", "1000101101111101", "1000111101111111", "1000011101111101", "1000011101111101", "1000101101111111", "1000011101111101", "1000011001111101", "1000001001111110", "1000011101111101", "1000011001111101", "1000011001111100", "1000100001111110", "1000101001111111", "1000111001111111", "1000110001111111", "1000110001111111", "1001001001111101", "1001011101111101", "1001101001111101", "1001110001111101", "1001110001111100", "1001110001111101", "1001111001111011", "1001111101111010", "1001111101111100", "1001111101111011", "1010000001111011", "1001111101111011", "1001111101111011", "1001110001111011", "1001101101111011", "1001100101111100", "1001011101111101", "1001010101111101", "1001010001111110", "1001001101111110", "1001000101111110", "1001000001111101", "1001000001111110", "1000111001111110", "1000110001111110", "1000101101111110", "1000110001111110", "1000111101111111", "1001001101111101", "1001000101111110", "1001000101111110", "1001010001111101", "1001001101111101", "1001000101111110", "1001110001111101", "1001100001111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100101111111", "1001111110000000", "1001111101111111", "1001111001111111", "1001111010000100", "1001100110000111", "1001100110000111", "1001011110000110", "1001100110000101", "1001110010000100", "1001110101111111", "1001011101111111", "1001010101111110", "1001101001111110", "1001101001111101", "1001100101111101", "1001101101111101", "1001110001111101", "1001100101111101", "1001100001111101", "1000101101111101", "1000101001111101", "1000100101111101", "1000100101111110", "1000110001111101", "1001000101111110", "1001001001111110", "1001000101111111", "1001100101111110", "1010000001111101", "1010000101111110", "1010000001111111", "1001111101111111", "1010000001111111", "1010000101111111", "1010001101111101", "1001101101111111", "1001010001111110", "1001001001111110", "1000100101111111", "1000011101111110", "1000010001111111", "1000010001111111", "1000011101111111", "1000000101111111", "1000100001111111", "1000011101111110", "1000010001111101", "1000010001111110", "1000011001111101", "1000010001111110", "1000001101111110", "1000000101111100", "1000000101111101", "1000000101111101", "0111111101111101", "1000001001111011", "1000001101111011", "1000011001111010", "1000010001111000", "1000010001111010", "1000011101111101", "1000101001111100", "1000101001111101", "1000100101111100", "1000110101111111", "1000011101111101", "1000010101111110", "1000101101111111", "1000011101111101", "1000011101111100", "1000001001111110", "1000011101111110", "1000011101111110", "1000011101111101", "1000100101111101", "1000110001111111", "1001000001111101", "1001000101111110", "1000101101111111", "1001001001111101", "1001011101111101", "1001101101111100", "1001101101111101", "1001110001111100", "1001111001111011", "1001111101111011", "1001111101111010", "1001111101111011", "1010000001111011", "1010000001111011", "1010000001111010", "1001111001111011", "1001110101111011", "1001101101111011", "1001101001111011", "1001100101111011", "1001011101111100", "1001010101111101", "1001010001111101", "1001001101111110", "1001000101111110", "1001000001111110", "1000111101111111", "1000110001111110", "1000101001111110", "1000100101111111", "1000110001111110", "1001001001111110", "1001000101111110", "1001000101111101", "1001001101111110", "1001001001111110", "1001001101111110", "1001110101111101", "1001100001111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001010101111111", "1001010001111111", "1001011001111111", "1001100101111111", "1001111110000000", "1010000110000000", "1010000110000000", "1001110010000110", "1001011110001000", "1001100010000111", "1001100010000110", "1001101010000100", "1001111010000001", "1001110101111111", "1001011001111111", "1001101001111110", "1001101101111101", "1001101101111101", "1001101101111101", "1001110001111101", "1001110001111101", "1001100101111101", "1001100101111101", "1000101101111111", "1000110001111101", "1000101001111101", "1000101001111101", "1000110001111101", "1000111101111101", "1001001101111110", "1001001001111110", "1001100101111110", "1010000001111110", "1010000101111110", "1001111101111111", "1001111101111111", "1001111101111111", "1010000001111111", "1010001101111101", "1001110101111101", "1001010001111101", "1000111001111111", "1000010001111101", "1000001001111111", "1000010001111110", "1000010001111111", "1000011101111111", "1000010101111110", "1000010001111111", "1000010001111110", "1000010101111110", "1000010001111101", "0111111101111111", "1000010001111110", "0111111101111111", "1000000101111101", "1000000101111110", "1000000101111101", "1000000101111101", "0111111101111101", "1000001101111011", "1000011001111001", "1000011101111001", "1000011001111010", "1000100001111010", "1000110101111101", "1000100101111011", "1000101001111110", "1000101101111110", "1000011101111101", "1000010101111110", "1000101101111111", "1000100001111110", "1000011001111101", "1000010001111101", "1000011101111110", "1000100001111110", "1000011101111101", "1000100101111111", "1000111001111111", "1001010001111101", "1001010101111101", "1000110001111111", "1001000101111110", "1001100001111101", "1001101001111101", "1001110001111100", "1001110101111100", "1001111101111010", "1010000001111010", "1010000001111011", "1010000001111100", "1001111101111011", "1001111101111011", "1010000001111011", "1001111101111011", "1001111001111011", "1001110001111011", "1001101101111010", "1001100101111011", "1001100101111011", "1001011101111100", "1001011001111101", "1001010101111101", "1001001001111110", "1001000101111110", "1000111101111110", "1000110001111101", "1000101001111110", "1000011101111110", "1000011101111110", "1000111001111110", "1001000101111110", "1001000101111110", "1001001001111101", "1001000101111110", "1001010101111110", "1001110101111110", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001010101111111", "1001011101111111", "1001101101111111", "1001111101111111", "1010000110000000", "1010000110000001", "1001100110000111", "1001011110001000", "1001011110000111", "1001100110000110", "1001110010000100", "1010000001111111", "1001110001111111", "1001100101111110", "1001110001111101", "1001110001111101", "1001110001111101", "1001110101111101", "1001110001111101", "1001101101111101", "1001100101111101", "1001100101111101", "1000100101111111", "1000101001111111", "1000101101111101", "1000100101111101", "1000101001111101", "1000111101111101", "1001000101111110", "1001000101111110", "1001100101111110", "1010000001111110", "1010000001111111", "1001111101111111", "1001111101111111", "1001111101111111", "1010000101111111", "1010001001111110", "1001110001111111", "1001010101111101", "1000110101111111", "1000001001111110", "0111111101111111", "1000001001111111", "1000010001111111", "0111111101111111", "1000010001111111", "1000001101111110", "1000010101111110", "1000010101111101", "1000011001111111", "1000001001111110", "1000010001111110", "1000000101111111", "1000000101111110", "1000010001111101", "1000001101111101", "1000001101111101", "1000000001111101", "0111111101111100", "1000010001111010", "1000100001111010", "1000001101111010", "1000010101111001", "1000111101111101", "1000011101111111", "1000101101111100", "1000100101111101", "1000011101111101", "1000011101111101", "1000101001111111", "1000100101111111", "1000011101111101", "1000010001111101", "1000011101111110", "1000100001111110", "1000011101111101", "1000100101111110", "1000111101111111", "1001011001111101", "1001011101111101", "1000111001111111", "1000111101111111", "1001011101111101", "1001110001111100", "1001111001111100", "1001111001111100", "1001111101111011", "1010000101111010", "1010000001111011", "1010000101111011", "1010000001111011", "1010000001111011", "1010000101111010", "1001111101111011", "1001111101111010", "1001110101111010", "1001101101111011", "1001101001111011", "1001100101111010", "1001100001111011", "1001011101111100", "1001010101111101", "1001010001111101", "1001001001111101", "1001000001111110", "1000111001111101", "1000101101111101", "1000011101111110", "1000011001111110", "1000011101111110", "1001000001111110", "1001001001111110", "1001000101111101", "1001000001111111", "1001011101111101", "1001101101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100101111111", "1001110101111111", "1010000101111111", "1010010010000001", "1001111110000101", "1001011110001000", "1001011110001000", "1001011110000111", "1001100110000101", "1001111010000010", "1001111101111111", "1001110001111110", "1001110001111101", "1001101101111101", "1001110001111101", "1001110101111101", "1001111001111101", "1001101101111101", "1001101001111101", "1001101001111101", "1001100001111110", "1000011101111111", "1000100101111111", "1000101001111110", "1000101101111101", "1000101101111101", "1000110101111101", "1001000001111110", "1001000101111110", "1001100101111110", "1010000101111101", "1010000101111110", "1001111001111111", "1001111101111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000001111110", "1001010001111111", "1000101101111111", "1000010001111101", "0111111101111111", "1000000101111111", "1000001101111111", "0111111101111111", "1000000001111111", "1000010001111110", "1000011101111101", "1000010001111101", "1000010101111110", "1000010001111101", "1000000101111111", "1000011101111110", "1000001101111110", "1000010001111101", "1000010001111101", "1000001101111100", "1000001001111010", "1000000001111100", "1000001001111011", "1000011101111010", "1000011001111001", "1000010101111001", "1000100101111101", "1000100101111110", "1000101001111011", "1000101001111101", "1000010101111110", "1000100101111101", "1000110001111111", "1000101101111110", "1000011101111101", "1000011001111101", "1000011101111110", "1000100001111110", "1000011101111101", "1000101101111110", "1001000001111110", "1001011101111101", "1001011101111101", "1000111101111111", "1001000001111101", "1001100001111100", "1001110101111100", "1001111001111100", "1001111101111011", "1010000101111010", "1010000101111011", "1010000101111011", "1010000101111100", "1010000001111100", "1010000001111011", "1010000101111010", "1010000001111010", "1001111101111010", "1001110101111011", "1001110001111010", "1001101101111010", "1001101001111011", "1001100001111100", "1001011101111100", "1001011001111101", "1001010001111101", "1001001001111101", "1000111101111101", "1000110001111110", "1000100101111110", "1000011101111111", "1000011001111111", "1000010001111111", "1000101101111110", "1001000101111110", "1001000101111111", "1000111101111111", "1001100101111101", "1001101101111110", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001101101111110", "1001111101111111", "1010010001111111", "1010000110000100", "1001110010000111", "1001011010001000", "1001011110001000", "1001100010000111", "1001110010000100", "1010000110000000", "1001111101111110", "1001110101111110", "1001110001111101", "1001110001111101", "1001110101111101", "1001111101111101", "1001110001111101", "1001100101111101", "1001101101111101", "1001100101111101", "1001011001111101", "1000011001111101", "1000011101111111", "1000101001111111", "1000110001111101", "1000101101111101", "1000110101111101", "1000111101111110", "1000111101111111", "1001100101111110", "1010000101111101", "1010000101111111", "1001111101111111", "1001111101111111", "1001111101111111", "1010000101111111", "1010001101111101", "1010000101111101", "1001011101111110", "1000100101111111", "1000010001111110", "0111111101111111", "1000001001111110", "1000000101111111", "0111111101111111", "1000000101111111", "1000001101111110", "1000011101111101", "1000010001111101", "1000010001111111", "1000010001111110", "1000010001111110", "1000001001111110", "1000010101111110", "1000010001111110", "1000010001111110", "1000001001111100", "1000001001111011", "1000000001111100", "1000000001111100", "1000011001111010", "1000010101111001", "1000011101111001", "1000011101111101", "1000110001111101", "1000101101111010", "1000100101111100", "1000010101111110", "1000100101111110", "1000110001111110", "1000110001111101", "1000100001111101", "1000011101111101", "1000100101111101", "1000100001111110", "1000100001111101", "1000110001111111", "1001001101111101", "1001011101111100", "1001011101111101", "1001000101111110", "1001000101111110", "1001100101111101", "1001111001111100", "1001111001111100", "1001111101111100", "1010000101111010", "1010000101111011", "1010000101111011", "1010000101111100", "1010000001111100", "1010000101111011", "1010000101111011", "1010000101111010", "1001111101111010", "1001111101111010", "1001111001111010", "1001110001111010", "1001101001111011", "1001101001111010", "1001100001111011", "1001011001111101", "1001010001111101", "1001001001111101", "1000111101111110", "1000110001111101", "1000100101111110", "1000011101111110", "1000011001111111", "1000010101111111", "1000011001111111", "1001000001111110", "1001000101111110", "1000111101111111", "1001110001111110", "1001101001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100101111111", "1001110001111111", "1010000101111111", "1010000010000100", "1001111110000100", "1001100110000111", "1001011010001001", "1001011110001000", "1001100110000110", "1001111110000100", "1010001001111111", "1001111101111110", "1001111001111101", "1001110101111101", "1001111001111101", "1001111101111101", "1001110101111101", "1001101001111101", "1001100101111101", "1001101101111101", "1001011101111101", "1001010101111101", "1000011101111100", "1000011101111111", "1000100101111111", "1000101101111101", "1000101101111101", "1000110001111101", "1000111101111110", "1000111101111111", "1001100101111110", "1010000101111110", "1010000101111110", "1001111101111111", "1001111101111111", "1001111101111111", "1010000001111111", "1010001101111110", "1010000101111101", "1001011001111101", "1000100101111111", "1000010101111110", "1000010101111110", "1000000101111111", "1000000101111111", "1000000001111111", "1000001001111110", "1000001101111110", "1000011101111011", "1000010101111101", "1000001001111110", "1000010001111111", "1000010101111110", "1000001101111110", "1000000101111111", "1000001001111110", "1000010001111101", "1000000101111101", "1000001101111011", "0111111101111100", "0111111101111101", "1000010001111010", "1000011101111001", "1000011001111010", "1000011101111010", "1000110001111110", "1000100101111010", "1000100001111100", "1000010101111101", "1000101101111110", "1000110101111110", "1000110001111110", "1000100101111110", "1000100001111110", "1000100101111110", "1000100001111110", "1000100101111111", "1000111101111111", "1001010101111101", "1001100101111100", "1001101001111100", "1001001001111101", "1001001001111101", "1001101001111101", "1001111001111100", "1001111101111100", "1010000101111010", "1010000101111010", "1010000101111010", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111010", "1010000101111010", "1010000001111011", "1001111101111010", "1001111001111011", "1001110001111011", "1001101101111010", "1001100101111010", "1001100001111011", "1001011101111011", "1001010101111101", "1001000101111101", "1000111101111101", "1000110001111101", "1000100101111101", "1000011101111110", "1000011001111110", "1000010101111111", "1000010001111111", "1000110001111111", "1001000001111110", "1001000001111110", "1001110101111110", "1001100101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001101001111111", "1001111101111111", "1001101110000101", "1001011110000110", "1001101110000101", "1001100110000111", "1001010110001000", "1001011110001000", "1001110010000110", "1010001110000001", "1010000101111111", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001100101111110", "1001011001111101", "1001010001111101", "1000100001111101", "1000011101111111", "1000100101111111", "1000101101111101", "1000101101111101", "1000110001111101", "1000111101111101", "1001000001111111", "1001100101111110", "1010000101111101", "1010000101111111", "1001111101111111", "1001111001111111", "1001111101111111", "1010000001111111", "1010001101111110", "1010000101111101", "1001010001111101", "1000100101111111", "1000011101111111", "1000001001111110", "0111111101111111", "1000000101111111", "1000000101111111", "1000000101111111", "1000011101111101", "1000100001111101", "1000010001111110", "0111111101111111", "1000010001111110", "1000010101111110", "1000001001111111", "1000000101111111", "1000010001111101", "1000001001111111", "1000001101111110", "1000001001111100", "1000001101111011", "1000000001111101", "1000010001111010", "1000011101111001", "1000011101111001", "1000110001111010", "1000100101111010", "1000011001111001", "1000010001111010", "1000011001111101", "1000110001111110", "1000110001111111", "1000110001111110", "1000100101111111", "1000101001111111", "1000100101111111", "1000100101111111", "1000110001111111", "1001010001111101", "1001101001111100", "1001101101111101", "1001101001111100", "1001000101111110", "1001010001111101", "1001110001111100", "1001111001111011", "1001111101111011", "1010000101111010", "1010000101111010", "1010000101111010", "1010000101111010", "1010000101111011", "1010000101111010", "1010000101111011", "1010000001111011", "1010000101111010", "1010000001111011", "1001111101111010", "1001111001111010", "1001110001111011", "1001110001111010", "1001101001111011", "1001100101111010", "1001011101111011", "1001010101111101", "1001001101111101", "1001000001111101", "1000110001111101", "1000100101111101", "1000011101111101", "1000011001111110", "1000011001111111", "1000010101111111", "1000011101111111", "1000111101111111", "1001000101111111", "1001111001111110", "1001011101111111", "1001011101111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100001111111", "1001110001111111", "1001111110000001", "1001011110000111", "1001011010000111", "1001100110000110", "1001011110000111", "1001011010001000", "1001100110000111", "1010000010000100", "1010010001111111", "1010001001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001111101111101", "1001111101111101", "1001110001111101", "1001110001111101", "1001101001111101", "1001011101111101", "1001010101111101", "1001010001111101", "1000011101111111", "1000011101111111", "1000100101111111", "1000101101111110", "1000101101111101", "1000110001111101", "1000111001111110", "1001000001111110", "1001100001111110", "1010000101111101", "1010000101111110", "1001111101111111", "1001111101111111", "1001111001111111", "1001111101111111", "1010000101111101", "1001111001111101", "1001001101111101", "1000101101111111", "1000010001111110", "1000001101111110", "1000000001111111", "1000000101111111", "1000001001111110", "1000010101111110", "1000010001111110", "1000011101111101", "1000010101111110", "1000000101111111", "1000010001111111", "1000010001111110", "1000000101111111", "1000000101111111", "1000010001111101", "1000000101111111", "1000010101111110", "1000000101111101", "1000001101111100", "1000001001111010", "1000011101111001", "1000100101111001", "1000100101111100", "1000011101111001", "1000011101111000", "1000101001111010", "1000100001111101", "1000110001111110", "1000111001111111", "1000110001111111", "1000101101111111", "1000101001111111", "1000101001111111", "1000101101111111", "1000101001111111", "1001000101111110", "1001011101111101", "1001110001111101", "1001110001111101", "1001101001111100", "1001000101111110", "1001011001111101", "1001110001111100", "1001111101111011", "1001111101111011", "1010000001111011", "1010000101111011", "1010000101111011", "1010000101111010", "1010000101111010", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111011", "1001111101111010", "1001111101111010", "1001110101111010", "1001110001111011", "1001101101111010", "1001101001111010", "1001100001111011", "1001010101111101", "1001010001111011", "1001000101111101", "1000110101111101", "1000101001111101", "1000100001111101", "1000011001111110", "1000011001111110", "1000010101111110", "1000010101111111", "1000111101111110", "1001001101111111", "1001111001111110", "1001011101111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001011101111111", "1001100101111111", "1001110101111111", "1001111110000001", "1001011110000111", "1001100110000111", "1001101110000111", "1001011010001000", "1001011110000111", "1001110110000111", "1010001110000001", "1010010001111110", "1010001101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001100101111101", "1001010101111101", "1001010101111101", "1001000101111110", "1000100001111111", "1000011101111111", "1000100001111111", "1000101001111110", "1000101101111101", "1000110001111101", "1000111001111110", "1000111101111111", "1001100001111110", "1010000101111101", "1010000101111110", "1001111101111111", "1001111101111111", "1001111001111111", "1001111101111111", "1010000101111101", "1001111101111101", "1001010001111101", "1000100101111110", "1000010101111101", "1000001001111110", "1000000101111111", "1000000101111110", "1000001101111111", "1000001101111110", "1000010001111101", "1000011101111111", "1000011001111111", "1000001001111110", "1000001001111111", "1000001101111111", "1000000101111111", "1000010001111101", "1000010001111110", "1000010001111110", "1000010001111110", "1000001001111110", "1000001001111110", "1000010001111010", "1000010001111010", "1000010101111010", "1000100101111100", "1000011101111110", "1000100101111110", "1000100101111110", "1000110001111101", "1000110001111101", "1000111101111101", "1001000101111101", "1000111101111101", "1000110001111111", "1000101001111111", "1000110001111111", "1000110001111111", "1001001101111101", "1001100001111101", "1001110001111100", "1001110001111100", "1001100101111101", "1001000101111110", "1001011101111101", "1001110101111100", "1001111101111011", "1010000001111011", "1010000101111011", "1010000101111011", "1010000101111010", "1010000101111011", "1010000101111010", "1010000101111010", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111010", "1010000101111010", "1001111101111010", "1001111001111010", "1001110101111010", "1001110001111010", "1001101001111010", "1001100001111011", "1001011101111100", "1001001101111101", "1001000101111101", "1000111101111101", "1000101101111101", "1000100101111101", "1000011101111101", "1000011001111110", "1000011001111110", "1000011001111110", "1000101101111111", "1001010101111110", "1001110101111111", "1001011101111111", "1001010101111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011001111111", "1001011101111111", "1001011101111111", "1001100101111111", "1001111001111111", "1001111110000010", "1001100110000111", "1001110010000111", "1001110010000111", "1001011010001000", "1001100010001000", "1001111110000101", "1010010101111111", "1010001101111110", "1010001001111101", "1001111101111101", "1001111001111101", "1001111101111101", "1001110101111101", "1001101101111101", "1001101001111101", "1001101001111101", "1001011101111101", "1001010101111101", "1001001101111101", "1001000101111110", "1000100001111111", "1000011001111111", "1000011101111111", "1000101001111110", "1000101001111110", "1000101101111101", "1000111001111101", "1000111101111111", "1001011101111110", "1010000101111101", "1010001001111110", "1001111101111111", "1001111001111111", "1001111001111111", "1001111101111111", "1010001001111110", "1001111101111101", "1001010001111101", "1000101101111111", "1000011101111111", "1000001101111101", "1000000101111111", "0111111101111111", "1000000001111111", "1000010101111101", "1000000101111111", "1000011001111110", "1000010101111101", "1000001101111110", "1000000101111111", "1000010001111110", "1000000101111111", "1000000101111111", "1000010001111110", "1000010001111101", "1000000101111111", "1000000101111101", "1000001101111101", "1000010001111011", "1000001101111010", "1000001001111011", "1000010001111010", "1000100001111011", "1000100101111110", "1000100001111101", "1000100001111110", "1000101101111110", "1000100101111111", "1000110001111111", "1000111001111111", "1000111101111111", "1000101101111111", "1000101001111111", "1000111101111111", "1001010101111101", "1001100101111100", "1001110001111100", "1001110001111101", "1001100101111101", "1001000101111110", "1001100101111101", "1001111001111100", "1001111101111100", "1010000001111011", "1010000101111010", "1010000101111011", "1010000101111010", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111100", "1010000101111011", "1010000101111010", "1010000101111010", "1001111101111010", "1001110101111010", "1001110001111011", "1001101001111010", "1001100101111010", "1001011101111100", "1001010001111100", "1001000101111101", "1000111101111101", "1000110001111101", "1000100101111101", "1000100001111101", "1000011001111110", "1000011001111110", "1000011001111110", "1000100001111110", "1001011101111110", "1001110001111111", "1001011001111111", "1001010101111111", "1001010101111111", "1001011001111111", "1001010101111111", "1001011001111111", "1001010101111111", "1001010101111111", "1001011001111111", "1001011001111111", "1001011101111111", "1001101001111111", "1001111101111111", "1010000110000000", "1001111110000110", "1001111110000111", "1001110010000111", "1001011010001000", "1001101010000111", "1010001110000010", "1010010001111110", "1010010001111101", "1010000101111101", "1001110101111101", "1001110001111101", "1001110101111101", "1001101001111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001011001111101", "1001010001111101", "1001001101111101", "1001000001111101", "1000011101111111", "1000011101111111", "1000100001111111", "1000101001111110", "1000101101111101", "1000101101111101", "1000110101111110", "1000111101111110", "1001011101111110", "1010000101111101", "1010000101111110", "1001111101111111", "1001111101111111", "1001111101111111", "1001111101111111", "1010001001111110", "1001111101111101", "1001011001111101", "1000110001111110", "1000011001111111", "1000000101111111", "1000001101111110", "1000001101111111", "1000100001111110", "1000010101111101", "1000000101111111", "1000010001111101", "1000010101111101", "1000001001111111", "1000000101111111", "1000000001111111", "1000000101111111", "1000010001111101", "1000001101111110", "1000010001111101", "1000010001111101", "1000010001111101", "1000000001111101", "0111111101111011", "1000000101111010", "1000001001111011", "1000001101111101", "1000010101111010", "1000100001111101", "1000100101111101", "1000010101111101", "1000110001111111", "1000100001111110", "1000110001111111", "1000100101111111", "1000101001111111", "1000100001111110", "1000101101111111", "1001001001111110", "1001011101111101", "1001100101111101", "1001110001111100", "1001110001111100", "1001011001111101", "1001010001111101", "1001110001111101", "1001111101111100", "1010000001111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111010", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111010", "1001111101111010", "1001111101111010", "1001110101111010", "1001101101111010", "1001100101111011", "1001100101111010", "1001010101111100", "1001001001111101", "1000111101111101", "1000110001111101", "1000100101111101", "1000100001111101", "1000011101111101", "1000011001111110", "1000011001111110", "1000011101111110", "1001100101111101", "1001110001111111", "1001011101111111", "1001011001111111", "1001011001111111", "1001010101111111", "1001010101111111", "1001010101111111", "1001010001111111", "1001010001111111", "1001011001111110", "1001011101111111", "1001011101111111", "1001101001111111", "1001111101111111", "1010001001111111", "1010001010000000", "1010000110000011", "1001101110000111", "1001011110001001", "1001110110000111", "1010010010000001", "1010010001111101", "1010000101111101", "1001111101111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001100001111101", "1001100101111101", "1001100101111101", "1001011101111101", "1001010101111101", "1001010001111101", "1001001001111101", "1001000001111101", "1000011101111111", "1000011101111101", "1000011101111111", "1000100101111111", "1000101001111110", "1000101101111101", "1000110001111110", "1000111101111110", "1001011101111110", "1010000101111101", "1010000101111110", "1001111101111111", "1001111101111111", "1001111001111111", "1001111101111111", "1010001101111101", "1001111001111101", "1001011101111101", "1000111101111110", "1000011101111110", "1000000101111111", "1000011101111111", "1000010001111111", "0111111101111111", "0111111101111111", "1000001001111110", "1000010101111110", "1000010001111101", "1000011001111101", "1000011101111110", "1000001001111111", "1000010101111110", "1000010001111111", "1000010001111110", "1000010001111101", "1000010001111110", "1000001101111101", "1000000101111111", "1000000101111101", "1000000101111100", "1000001001111011", "1000010001111110", "1000001101111101", "1000010001111010", "1000010001111010", "1000011101111110", "1000100101111111", "1000011101111110", "1000100101111111", "1000100001111111", "1000011101111110", "1000100101111110", "1000111001111111", "1001010001111101", "1001100101111100", "1001101101111100", "1001110001111100", "1001101001111100", "1001000101111110", "1001011101111101", "1001111001111011", "1010000001111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111010", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111010", "1010000001111010", "1001111101111010", "1001110101111010", "1001110001111010", "1001101001111010", "1001100101111010", "1001011101111100", "1001001101111101", "1001000001111101", "1000110001111101", "1000101001111101", "1000100001111101", "1000011101111110", "1000011101111101", "1000011001111110", "1000011101111101", "1001010101111101", "1001101101111111", "1001011001111111", "1001010101111111", "1001010101111111", "1001011001111111", "1001011001111111", "1001010101111111", "1001010101111111", "1001010101111111", "1001010101111111", "1001011001111111", "1001100001111111", "1001110001111111", "1001111101111111", "1010001001111110", "1010001001111111", "1010000010000001", "1001101010001000", "1001100010001001", "1010000010000110", "1010010101111111", "1010010001111101", "1010000001111101", "1001110101111101", "1001110001111101", "1001101101111101", "1001011101111101", "1001011101111101", "1001100101111101", "1001011101111101", "1001010101111101", "1001010001111101", "1001001101111101", "1001000101111101", "1000111001111110", "1000011101111111", "1000011001111101", "1000011101111111", "1000100101111110", "1000101101111101", "1000110001111101", "1000110101111101", "1000111101111110", "1001011101111110", "1010000001111101", "1010000101111101", "1001111101111111", "1001111101111111", "1001111101111111", "1010000001111111", "1010001001111110", "1001111101111101", "1001010101111101", "1000111101111110", "1000011001111110", "1000001001111110", "1000001101111110", "0111111101111111", "0111111101111111", "1000000001111111", "1000010001111110", "1000010101111101", "1000001001111110", "1000011101111110", "1000000101111111", "1000010001111110", "1000001101111110", "0111111101111111", "1000010001111110", "1000010001111110", "1000010001111110", "1000001001111011", "1000001101111101", "1000010101111101", "1000001101111110", "1000010001111101", "1000010101111110", "1000011101111100", "1000100001111101", "1000100001111101", "1000101001111111", "1000011101111110", "1000011101111110", "1000011101111101", "1000011101111101", "1000011101111101", "1000101101111111", "1001000001111111", "1001011001111101", "1001100101111100", "1001101101111100", "1001101101111100", "1001011101111101", "1001000001111110", "1001101001111100", "1001111101111100", "1010000001111011", "1010000101111010", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111010", "1010000001111010", "1010000001111010", "1001111001111010", "1001110101111010", "1001101101111010", "1001101001111010", "1001011101111011", "1001010001111101", "1001001001111100", "1000111101111101", "1000101101111101", "1000100001111101", "1000011101111110", "1000011001111110", "1000011101111110", "1000011101111101", "1000111101111101", "1001100101111111", "1001011001111111", "1001010101111111", "1001010101111110", "1001010101111111", "1001010101111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001010001111111", "1001011001111111", "1001100001111111", "1001110001111111", "1001111101111111", "1010000001111111", "1010000101111111", "1001111110000100", "1001100110001000", "1001101110001000", "1010001010000010", "1010010101111101", "1010000101111101", "1001110001111101", "1001101101111101", "1001101101111101", "1001011101111101", "1001011101111101", "1001100101111101", "1001011101111101", "1001011001111101", "1001010101111101", "1001010001111101", "1001001001111101", "1000111101111110", "1000110001111111", "1000011101111111", "1000011101111100", "1000011101111111", "1000100101111111", "1000110001111101", "1000101101111101", "1000110001111101", "1000111101111110", "1001011001111110", "1001111101111101", "1010000101111101", "1001111101111111", "1001111001111111", "1001111001111111", "1001111101111111", "1010001001111110", "1010000101111101", "1001011001111101", "1001000001111101", "1000010001111110", "1000011001111101", "1000001101111110", "0111111101111111", "0111111101111111", "1000010001111111", "1000001001111111", "1000001101111111", "1000001101111110", "1000011101111110", "1000010001111101", "1000000101111111", "1000001001111110", "1000001101111110", "1000001101111111", "1000001101111110", "1000010001111100", "1000010001111011", "1000001001111010", "1000010001111110", "1000010101111110", "1000011101111110", "1000100001111110", "1000100101111101", "1000100101111110", "1000100101111101", "1000100101111111", "1000010001111110", "1000011101111101", "1000010101111101", "1000011001111101", "1000100101111101", "1000111101111111", "1001001101111110", "1001100001111100", "1001101001111100", "1001101001111100", "1001100101111100", "1000111101111110", "1001010001111101", "1001110001111101", "1001111101111101", "1001111101111100", "1010000101111010", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111100", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111011", "1010000001111010", "1001111101111010", "1001110101111010", "1001110001111010", "1001101001111011", "1001100101111010", "1001011001111100", "1001001101111100", "1000111101111101", "1000110001111101", "1000100101111101", "1000100001111101", "1000011001111110", "1000011001111110", "1000011101111101", "1000100101111101", "1001011101111110", "1001011101111111", "1001011001111101", "1001010101111101", "1001010001111110", "1001010001111111", "1001010001111110", "1001001101111110", "1001001001111111", "1001001001111111", "1001010001111111", "1001100001111111", "1001110101111111", "1001111110000000", "1010000010000001", "1010000110000001", "1001110110000110", "1001011110001000", "1001111010000110", "1010010001111111", "1010000101111101", "1001110001111101", "1001100101111101", "1001100101111101", "1001100101111101", "1001011101111101", "1001100001111101", "1001011101111101", "1001010101111101", "1001010101111101", "1001010101111101", "1001010001111101", "1001000101111101", "1000111001111110", "1000101101111111", "1000101001111111", "1000011101111111", "1000100001111111", "1000101001111111", "1000110001111101", "1000110001111101", "1000110101111101", "1000111101111101", "1001010101111110", "1001111101111111", "1010000101111110", "1001111101111111", "1001111001111111", "1001111001111111", "1001111101111111", "1010000101111110", "1001111101111101", "1001011001111101", "1001000001111101", "1000010101111101", "1000010101111110", "1000000101111111", "0111111101111111", "1000010001111111", "1000010001111110", "1000000101111111", "1000001101111110", "1000010001111110", "1000011001111111", "1000011001111101", "1000010001111101", "1000001101111110", "1000010001111110", "1000010001111101", "1000000101111111", "1000010001111101", "1000001101111101", "1000010001111010", "1000000101111010", "1000011101111101", "1000100101111101", "1000100101111101", "1000011101111111", "1000010101111101", "1000100001111110", "1000010101111101", "1000011001111101", "1000010001111101", "1000010101111101", "1000011001111101", "1000101101111111", "1001000101111110", "1001011001111101", "1001100101111101", "1001101001111100", "1001101001111100", "1001001101111110", "1000111101111111", "1001100101111101", "1001111001111101", "1010000001111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111010", "1010000001111010", "1001111101111010", "1001110101111010", "1001101101111010", "1001100101111011", "1001011101111100", "1001010001111100", "1001000101111101", "1000110101111101", "1000101001111101", "1000100101111101", "1000011101111101", "1000011001111110", "1000011001111110", "1000011101111101", "1001010001111101", "1001011101111111", "1001011101111111", "1001011101111110", "1001011001111101", "1001010001111110", "1001000101111111", "1001000001111111", "1000111101111111", "1000110001111111", "1000111101111111", "1001010101111111", "1001110001111111", "1001111110000100", "1010000010000100", "1010000110000011", "1001110010000111", "1001101110000111", "1010000110000011", "1010001001111110", "1001110001111101", "1001011101111101", "1001100001111101", "1001011101111101", "1001011001111101", "1001011101111101", "1001011101111101", "1001011001111101", "1001010001111101", "1001010001111101", "1001010001111101", "1001001001111101", "1000111101111101", "1000110001111111", "1000101001111111", "1000111001111111", "1000110101111111", "1000111101111110", "1000111001111110", "1000110101111101", "1000110001111101", "1000110001111101", "1000111001111110", "1001010101111110", "1001111101111101", "1010000001111110", "1001111101111111", "1001111001111111", "1001111001111111", "1001111101111111", "1010000101111111", "1001110001111110", "1001011101111101", "1000110001111110", "1000011101111110", "1000001101111111", "1000001001111110", "1000001101111111", "1000001001111111", "1000010001111110", "1000000101111111", "1000010001111110", "1000010101111110", "1000011001111101", "1000011001111101", "1000010001111110", "1000010001111101", "1000000101111111", "1000010001111110", "1000010001111110", "1000010101111110", "1000010001111110", "1000011001111100", "1000000101111010", "1000001001111010", "1000011001111101", "1000110001111101", "1000100101111101", "1000011101111101", "1000011101111110", "1000010001111101", "1000010001111101", "1000010001111101", "1000010001111101", "1000011101111101", "1000111101111111", "1001010001111101", "1001100001111100", "1001100101111101", "1001100101111100", "1001011101111101", "1000110001111111", "1001010101111101", "1001110101111101", "1001111101111100", "1010000101111010", "1010000101111011", "1010000101111010", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111010", "1010000101111010", "1010000001111010", "1001111101111010", "1001110001111011", "1001101101111010", "1001100101111011", "1001011001111100", "1001001001111101", "1000111101111101", "1000110001111100", "1000100101111100", "1000011101111101", "1000011101111101", "1000011101111101", "1000100001111101", "1000111101111101", "1001011001111101", "1001011101111110", "1001011101111111", "1001011001111111", "1001010101111101", "1001010001111110", "1001000101111110", "1000111101111111", "1000101101111111", "1000101001111111", "1001000001111111", "1001111010000010", "1001111110000111", "1010000110000101", "1010000110000011", "1001110110000111", "1001111110000110", "1010001001111111", "1001110001111110", "1001011101111101", "1001011001111101", "1001011101111101", "1001010101111101", "1001011001111101", "1001011001111101", "1001010001111101", "1001010001111101", "1001001101111110", "1001010001111101", "1001010001111101", "1001000101111101", "1000111001111110", "1000110001111111", "1000101001111111", "1001000001111110", "1001001001111101", "1001001001111101", "1001000001111101", "1000110101111101", "1000101101111110", "1000101101111111", "1000111001111101", "1001010001111110", "1001111101111110", "1010000001111101", "1001111101111111", "1001111101111111", "1001111101111111", "1001111101111111", "1010000101111110", "1001110001111101", "1001011101111101", "1000110001111110", "1000011101111110", "1000010101111101", "1000010001111111", "0111111101111111", "1000000001111111", "1000000101111111", "0111111101111111", "1000000101111111", "1000010101111110", "1000010001111110", "1000011001111101", "1000010001111110", "1000000101111111", "1000000101111111", "1000001001111110", "1000010101111111", "1000011001111110", "1000011001111110", "1000011001111110", "1000011101111101", "1000010001111010", "1000011001111010", "1000011101111101", "1000100101111100", "1000100001111101", "1000010001111101", "1000010001111101", "1000001101111110", "1000000101111111", "1000011101111101", "1000110001111111", "1001000101111110", "1001011101111101", "1001100101111101", "1001100101111101", "1001011101111101", "1000110001111111", "1001001001111101", "1001110001111100", "1001111101111100", "1001111101111100", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111100", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010001001111010", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111100", "1010000101111011", "1010000101111010", "1010000001111010", "1001111101111010", "1001110001111011", "1001101101111011", "1001100101111011", "1001011101111100", "1001010001111101", "1001000001111101", "1000110001111101", "1000100101111101", "1000100001111101", "1000100001111100", "1000011101111101", "1000100101111101", "1000101101111101", "1001010101111101", "1001011001111101", "1001011101111110", "1001011101111111", "1001011001111111", "1001010101111101", "1001001101111110", "1001000101111110", "1000111101111111", "1000111001111111", "1001001001111111", "1010000110000001", "1010000110000111", "1010000110000101", "1010000110000100", "1010000110000100", "1010000101111111", "1001110001111110", "1001010101111110", "1001010001111110", "1001010101111101", "1001010101111101", "1001010101111101", "1001011001111101", "1001010001111101", "1001001001111101", "1001001001111101", "1001001101111101", "1001010001111101", "1001001101111101", "1001000001111110", "1000111001111110", "1000110001111111", "1000101101111111", "1000111001111111", "1001001001111101", "1001001101111101", "1001000101111101", "1000110101111101", "1000101101111110", "1000101101111110", "1000111001111101", "1001010001111110", "1001111001111110", "1010000001111110", "1001111101111111", "1001111001111111", "1001111001111111", "1001111101111111", "1010000101111111", "1001101101111101", "1001011101111101", "1000101101111101", "1000010101111110", "1000000101111111", "0111111101111111", "0111111101111111", "1000000101111111", "1000010001111110", "1000000101111111", "1000000001111111", "1000000101111111", "1000010101111101", "1000010001111101", "1000011001111110", "1000001101111110", "1000001001111110", "1000010101111101", "1000010001111110", "1000011101111111", "1000010101111110", "1000011101111101", "1000011101111110", "1000100001111101", "1000011001111101", "1000011001111100", "1000011101111110", "1000010101111101", "1000001101111110", "1000001001111110", "1000000101111111", "1000010001111101", "1000100101111110", "1001000001111111", "1001010001111101", "1001011101111101", "1001100101111100", "1001001101111101", "1000101001111111", "1001001001111101", "1001100101111101", "1001111001111100", "1001111101111100", "1001111101111100", "1010000101111011", "1010000101111010", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111010", "1010000001111010", "1001110101111010", "1001110001111010", "1001101001111100", "1001100101111011", "1001011001111100", "1001001001111100", "1000111101111100", "1000101101111101", "1000100101111101", "1000011101111101", "1000011101111101", "1000100001111101", "1000100101111101", "1001001001111101", "1001010101111101", "1001010101111110", "1001011001111110", "1001011001111111", "1001010101111111", "1001010001111110", "1001001001111111", "1001001001111110", "1001001101111110", "1001011101111110", "1001111101111111", "1001111010000110", "1001111110000111", "1010001010000010", "1010000101111111", "1001101101111110", "1001010101111110", "1001010001111110", "1001010101111101", "1001010001111101", "1001010001111101", "1001011001111101", "1001010001111101", "1001000101111101", "1001000101111101", "1001001001111101", "1001010001111101", "1001010001111101", "1001000101111101", "1001000001111101", "1000110101111110", "1000101101111111", "1000101101111111", "1000100101111111", "1001000001111110", "1001000101111101", "1001000001111101", "1000110001111101", "1000110001111101", "1000101101111110", "1000111001111110", "1001010001111110", "1001111001111110", "1010000101111101", "1001111101111111", "1001111001111111", "1001111001111111", "1001111101111111", "1010000101111110", "1001101001111110", "1001011101111101", "1000100001111101", "1000010001111110", "1000001001111110", "1000001001111110", "1000010001111101", "1000001001111110", "1000010101111110", "1000001001111110", "1000000101111111", "1000011001111110", "1000011001111101", "1000010101111101", "1000011001111111", "1000010001111110", "1000010001111110", "1000011001111110", "1000011001111110", "1000011001111110", "1000011001111101", "1000010101111110", "1000011001111110", "1000011101111100", "1000011101111101", "1000011001111111", "1000011001111101", "1000000101111111", "1000010001111110", "1000000001111111", "1000000101111111", "1000011101111101", "1000110101111111", "1001001001111110", "1001010001111101", "1001000001111110", "1000110001111110", "1000111001111101", "1001011001111101", "1001101001111100", "1001110001111100", "1001111001111101", "1001111101111100", "1010000001111011", "1010000101111011", "1010000101111011", "1010001001111010", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111011", "1010000101111100", "1010000101111100", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000001111010", "1001111001111010", "1001110101111010", "1001101101111011", "1001100101111011", "1001011101111100", "1001010001111100", "1000111101111100", "1000110101111101", "1000101001111100", "1000011101111101", "1000011101111101", "1000011101111101", "1000100101111100", "1001000001111101", "1001010001111110", "1001010001111110", "1001010101111101", "1001011001111110", "1001010001111111", "1001010001111110", "1001010001111110", "1001010001111110", "1001011101111110", "1001101101111110", "1001111101111111", "1001110010000011", "1001111110000001", "1001111101111111", "1001100101111110", "1001011001111101", "1001010001111110", "1001010101111101", "1001010001111101", "1001010101111101", "1001010101111101", "1001010001111101", "1001000101111101", "1001000001111110", "1001000101111101", "1001001101111101", "1001010001111110", "1001001101111101", "1001000101111101", "1000111101111101", "1000110001111111", "1000101101111111", "1000101001111111", "1000100001111111", "1000110001111111", "1000111101111110", "1000111001111101", "1000110001111101", "1000101101111110", "1000101101111110", "1000111001111101", "1001010001111110", "1001110101111110", "1010000101111110", "1001111101111111", "1001111001111111", "1001111001111111", "1001111101111111", "1010000101111110", "1001110001111101", "1001001001111101", "1000011101111101", "1000010001111101", "1000001001111110", "1000001101111110", "1000011001111110", "1000010001111101", "1000010001111110", "1000010001111110", "1000010001111101", "1000011101111111", "1000011001111101", "1000010101111110", "1000011101111110", "1000011101111101", "1000010001111110", "1000010001111110", "1000011001111110", "1000001101111111", "1000011001111101", "1000011001111110", "1000010001111101", "1000011101111011", "1000011101111010", "1000100001111110", "1000010001111110", "1000000101111111", "1000000101111111", "1000000001111111", "1000010001111101", "1000011101111101", "1000100101111110", "1000100101111101", "1000110001111101", "1000111101111101", "1001010101111101", "1001100101111101", "1001110001111100", "1001111001111100", "1001111001111100", "1001111101111011", "1001111101111100", "1010000001111011", "1010000101111011", "1010000101111010", "1010001001111010", "1010000101111011", "1010001001111010", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010001001111011", "1010001001111010", "1010001001111010", "1010001001111010", "1010000101111011", "1010000001111011", "1001111101111010", "1001110101111011", "1001110001111011", "1001100101111011", "1001100001111011", "1001010101111101", "1001001001111100", "1000111101111101", "1000101101111101", "1000100101111101", "1000011101111110", "1000011101111101", "1000100001111101", "1000110101111101", "1001001101111111", "1001010001111110", "1001010001111110", "1001010001111110", "1001010001111110", "1001010001111110", "1001010001111111", "1001011001111111", "1001101001111110", "1001110101111110", "1001111101111110", "1010000101111110", "1001111001111110", "1001101001111101", "1001100001111101", "1001011101111101", "1001011101111101", "1001010101111101", "1001010001111101", "1001010101111101", "1001010001111101", "1001000101111101", "1001000001111110", "1000111101111110", "1001001001111101", "1001010101111101", "1001010001111101", "1001000101111101", "1001000001111101", "1000110101111110", "1000101101111111", "1000101101111111", "1000100101111111", "1000100001111111", "1000101001111111", "1000110101111101", "1000110001111101", "1000110001111101", "1000101101111110", "1000101101111110", "1000111001111101", "1001010001111110", "1001110101111110", "1010000101111101", "1001111101111111", "1001111001111111", "1001111101111111", "1001111101111111", "1010000101111111", "1001110001111101", "1000111001111111", "1000011101111111", "1000010101111101", "1000001101111110", "1000001101111110", "1000011101111101", "1000010001111101", "1000010101111110", "1000001101111101", "1000010001111101", "1000011001111110", "1000011001111110", "1000010101111101", "1000011101111101", "1000011101111100", "1000011001111101", "1000001101111110", "1000100101111101", "1000001101111110", "1000010101111111", "1000100001111101", "1000011001111110", "1000011101111100", "1000011101111101", "1000011101111101", "1000010101111101", "1000000101111111", "1000000001111111", "1000001001111110", "1000011101111101", "1000101001111101", "1000111101111110", "1001010001111101", "1001011101111101", "1001100101111101", "1001110001111100", "1001110001111100", "1001111001111100", "1001111001111100", "1001111101111100", "1001111101111100", "1001111101111100", "1010000001111011", "1010000101111011", "1010001101111010", "1010001101111010", "1010001001111010", "1010000101111100", "1010001001111010", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010001001111010", "1010001001111010", "1010000101111011", "1010000101111011", "1010000101111010", "1001111101111010", "1001111101111010", "1001110001111010", "1001101101111010", "1001100001111011", "1001011001111100", "1001001101111100", "1001000101111100", "1000110001111101", "1000101001111101", "1000100001111101", "1000011101111101", "1000100001111101", "1000101001111101", "1001001101111101", "1001001101111110", "1001010001111110", "1001010001111110", "1001010001111110", "1001010001111110", "1001010101111110", "1001100001111110", "1001110001111110", "1001111101111101", "1001111101111101", "1001110101111101", "1001110001111101", "1001110001111101", "1001110001111101", "1001101101111101", "1001100001111101", "1001011001111101", "1001010101111101", "1001010001111101", "1001000101111101", "1001000101111101", "1001000101111101", "1001000101111101", "1001010001111101", "1001010001111110", "1001001001111101", "1001000101111101", "1000111101111101", "1000110001111110", "1000101101111111", "1000101001111111", "1000100101111111", "1000100001111111", "1000100101111111", "1000101101111111", "1000110001111101", "1000110001111110", "1000110001111110", "1000101101111111", "1000111001111111", "1001010001111110", "1001110001111110", "1010000101111110", "1001111101111111", "1001111101111111", "1001111001111111", "1001111101111111", "1010000001111110", "1001011001111101", "1000110101111110", "1000011101111111", "1000010101111101", "1000010001111101", "1000010001111101", "1000011001111101", "1000011001111101", "1000010101111110", "1000010001111101", "1000010001111101", "1000011001111101", "1000010101111101", "1000010001111101", "1000011101111100", "1000011001111101", "1000011001111011", "1000010001111110", "1000011101111101", "1000011101111110", "1000001001111111", "1000101001111110", "1000011101111101", "1000011001111110", "1000011101111100", "1000010101111101", "1000001101111111", "1000000101111111", "1000010001111101", "1000011101111101", "1000101001111111", "1001000101111110", "1001010101111101", "1001100001111101", "1001101101111101", "1001101101111101", "1001110001111100", "1001111001111100", "1001111101111100", "1001111101111100", "1001111101111101", "1001111101111101", "1001111101111100", "1010000101111011", "1010000101111011", "1010001101111010", "1010001001111010", "1010001001111010", "1010001001111010", "1010001101111010", "1010001001111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000001111010", "1001111101111010", "1001110001111011", "1001101101111010", "1001100101111011", "1001011101111011", "1001010001111100", "1001000101111101", "1000111101111101", "1000110001111101", "1000100101111100", "1000100101111100", "1000100101111101", "1000100101111101", "1001000101111101", "1001001001111110", "1001001101111111", "1001010001111110", "1001010001111110", "1001010001111110", "1001011101111101", "1001101001111110", "1001111001111110", "1010000001111101", "1001111101111101", "1001111101111101", "1001111001111101", "1001111001111101", "1001111101111101", "1001110001111101", "1001100001111101", "1001011001111101", "1001010001111101", "1001000101111101", "1001000001111110", "1001000001111110", "1001000101111110", "1001010001111101", "1001010101111101", "1001010001111101", "1001000101111101", "1000111101111101", "1000111001111110", "1000101101111111", "1000101001111111", "1000101001111111", "1000110001111111", "1000011101111111", "1000100101111111", "1000101001111111", "1000101001111110", "1000110101111110", "1000110001111111", "1000101001111111", "1000110001111111", "1001001101111111", "1001110001111110", "1010000101111110", "1001111101111111", "1001111101111111", "1001111101111111", "1001111101111111", "1010000001111101", "1001011101111100", "1000110101111111", "1000100101111111", "1000011101111110", "1000001101111110", "1000010101111101", "1000011101111110", "1000011101111111", "1000011001111111", "1000010001111101", "1000010101111101", "1000010101111101", "1000011101111110", "1000011001111110", "1000100101111101", "1000100101111101", "1000011101111011", "1000011101111101", "1000011001111110", "1000011101111101", "1000010101111110", "1000100101111110", "1000101001111101", "1000011101111110", "1000100101111110", "1000010001111101", "1000011001111101", "1000001001111110", "1000011101111101", "1000101101111111", "1001000101111110", "1001010101111101", "1001100001111101", "1001101001111100", "1001110001111100", "1001110001111100", "1001110101111100", "1001111101111100", "1001111101111100", "1001111101111100", "1001111101111100", "1001111101111011", "1010000101111011", "1010000101111100", "1010001001111010", "1010001101111010", "1010001101111010", "1010001001111010", "1010001001111010", "1010001101111011", "1010001101111010", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010000001111010", "1010000001111010", "1001111001111010", "1001110001111011", "1001101101111011", "1001100101111100", "1001100001111011", "1001011001111011", "1001001001111100", "1001000001111100", "1000110001111101", "1000101001111100", "1000100101111101", "1000100001111101", "1000100101111101", "1000111101111101", "1001000101111110", "1001001001111110", "1001010001111110", "1001001101111110", "1001011001111101", "1001100101111110", "1001110101111101", "1010000101111101", "1010001001111101", "1010000101111101", "1010000101111101", "1010001001111101", "1010010001111100", "1001111101111101", "1001101101111101", "1001100001111101", "1001010001111101", "1001000101111101", "1001000101111110", "1001000101111101", "1001000101111110", "1001001101111101", "1001011001111101", "1001010101111101", "1001001101111101", "1001000001111101", "1000110101111101", "1000101101111111", "1000101001111111", "1000101001111111", "1000110001111111", "1001000001111110", "1000100101111111", "1000100101111111", "1000101001111111", "1000101001111110", "1000111001111110", "1000110001111111", "1000101101111111", "1000110001111111", "1001001101111111", "1001110001111110", "1010000101111110", "1001111101111111", "1001111101111111", "1001111001111111", "1001111101111111", "1001111101111110", "1001011001111101", "1000110001111111", "1000100001111111", "1000011101111111", "1000010001111111", "1000011101111110", "1000100001111111", "1000100101111111", "1000100001111111", "1000011101111111", "1000011101111111", "1000011101111100", "1000011101111111", "1000100101111110", "1000101001111101", "1000100101111101", "1000100101111101", "1000011101111100", "1000011101111110", "1000100101111100", "1000011101111111", "1000011001111111", "1000101101111110", "1000011101111110", "1000011101111110", "1000011101111110", "1000100101111100", "1000100101111101", "1000110001111111", "1001000101111110", "1001010001111101", "1001011101111101", "1001100101111100", "1001110001111100", "1001110001111100", "1001110101111100", "1001111001111100", "1001111101111100", "1001111101111100", "1001111101111101", "1001111101111100", "1001111101111100", "1010000101111100", "1010000101111100", "1010001001111010", "1010001101111010", "1010001101111010", "1010001101111010", "1010001001111010", "1010010001111010", "1010001001111010", "1010001001111011", "1010000101111100", "1010000101111011", "1010000101111011", "1010001001111010", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111010", "1010000101111011", "1010000101111010", "1010000001111010", "1010000001111010", "1001111101111010", "1001110001111011", "1001110001111010", "1001101001111011", "1001100101111011", "1001011001111100", "1001010001111011", "1001000001111100", "1000111001111100", "1000110001111100", "1000101001111100", "1000100101111101", "1000100101111101", "1000110001111101", "1001010101111100", "1001001001111110", "1001001101111111", "1001010001111101", "1001100001111101", "1001101101111110", "1001111101111110", "1010010001111101", "1010010001111100", "1010010001111101", "1010010101111101", "1010010101111101", "1010010001111101", "1001111001111101", "1001101001111101", "1001011001111101", "1001000101111110", "1001000101111101", "1001001001111101", "1001000101111101", "1001001101111101", "1001011001111101", "1001011001111101", "1001010101111100", "1001000101111101", "1000111001111110", "1000101101111111", "1000101001111111", "1000101001111111", "1000101101111111", "1001000101111101", "1001011001111101", "1000101001111111", "1000100101111111", "1000101101111111", "1000101001111111", "1000110001111111", "1000110001111111", "1000101001111111", "1000110001111111", "1001001001111110", "1001110001111110", "1010000101111101", "1001111101111111", "1001111001111111", "1001111001111111", "1001111001111111", "1001111101111110", "1001010001111101", "1000111001111110", "1000011101111111", "1000100101111111", "1000010101111110", "1000011101111110", "1000100101111111", "1000101001111111", "1000100101111111", "1000100101111110", "1000100101111101", "1000100101111100", "1000011101111111", "1000100001111110", "1000101101111101", "1000100001111101", "1000101101111110", "1000100101111101", "1000100101111101", "1000100001111100", "1000010101111110", "1000011001111110", "1000100101111110", "1000100101111111", "1000100101111110", "1000100001111110", "1000011101111110", "1000110001111111", "1001000001111110", "1001010001111101", "1001010101111101", "1001100001111100", "1001101001111100", "1001110001111100", "1001110001111100", "1001111001111100", "1001111001111101", "1001111101111101", "1001111101111100", "1001111101111101", "1001111101111100", "1010000001111100", "1010000101111011", "1010000101111011", "1010001001111010", "1010001101111010", "1010001101111010", "1010001101111010", "1010001101111010", "1010001101111010", "1010001101111010", "1010001001111011", "1010001001111011", "1010000101111100", "1010001001111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111011", "1010000101111010", "1010000101111010", "1001111101111010", "1001111001111010", "1001111001111011", "1001110101111010", "1001101101111010", "1001101101111010", "1001100101111010", "1001011101111011", "1001001101111100", "1001000101111100", "1000111101111100", "1000110001111100", "1000100101111101", "1000100101111101", "1000100101111101", "1000101101111101", "1001110001110110", "1001110001110111", "1001011101111100", "1001010101111110", "1001100101111110", "1001111001111101", "1010001101111101", "1010010101111101", "1010010001111101", "1010010101111101", "1010010101111110", "1010010101111101", "1010000101111101", "1001110001111101", "1001011101111101", "1001000101111101", "1001000101111110", "1001000101111101", "1001001001111101", "1001010001111101", "1001011001111101", "1001011101111101", "1001010101111101", "1001001101111101", "1000111101111101", "1000101101111111", "1000101001111111", "1000100101111111", "1000101001111111", "1001000001111110", "1001010101111101", "1001011101111101", "1000110001111111", "1000101101111111", "1000110001111111", "1000110001111111", "1000110001111110", "1000101001111101", "1000101001111111", "1000110001111110", "1001001101111101", "1001110101111101", "1010000101111110", "1001111101111111", "1001111001111111", "1001111001111111", "1001111001111111", "1010000001111110", "1001010001111101", "1000111101111111", "1000100101111111", "1000101001111111", "1000101001111110", "1000100101111110", "1000100101111111", "1000100101111111", "1000100001111111", "1000100101111111", "1000100101111110", "1000011101111101", "1000010101111101", "1000011101111110", "1000101101111101", "1000011101111101", "1000101101111110", "1000110001111101", "1000100001111101", "1000101001111100", "1000011101111101", "1000010001111110", "1000011101111110", "1000100101111111", "1000011101111110", "1000010101111110", "1000100001111110", "1000111101111111", "1001001101111101", "1001011001111101", "1001011101111101", "1001100101111100", "1001101101111100", "1001110101111011", "1001111001111100", "1001111101111100", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1001111101111101", "1010000101111011", "1010000101111011", "1010001001111010", "1010001101111010", "1010001001111010", "1010001101111010", "1010001101111010", "1010001001111011", "1010001001111010", "1010001101111010", "1010001101111011", "1010001101111011", "1010001101111010", "1010001101111011", "1010000101111011", "1010000101111011", "1010001001111010", "1010001001111010", "1010000101111011", "1010000101111011", "1010000101111010", "1010000101111010", "1010000001111010", "1001111101111010", "1001110101111011", "1001110101111011", "1001110001111010", "1001101101111011", "1001101001111011", "1001011101111011", "1001011101111011", "1001010001111100", "1001000101111101", "1000111101111100", "1000110101111100", "1000101101111101", "1000100101111100", "1000100101111101", "1000101001111101", "1001001101111100", "1001100101111010", "1001110001110110", "1001110101110111", "1001111101111010", "1010001001111100", "1010010101111100", "1010010101111101", "1010010101111101", "1010010101111110", "1010010101111110", "1010001001111101", "1001111001111101", "1001100001111101", "1001001101111110", "1001001001111101", "1001001101111101", "1001010001111101", "1001010101111101", "1001011101111101", "1001100101111101", "1001011101111101", "1001001001111101", "1000111101111101", "1000110001111111", "1000100101111111", "1000100101111111", "1000101001111111", "1000111101111101", "1001010001111101", "1001011101111100", "1001100101111100"
	);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			data <= rom(to_integer(unsigned(address)));
		end if;
	end process;
end Behavioral;